CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
10 10 30 70 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
42
13 Logic Switch~
5 63 353 0 10 11
0 35 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 64 294 0 10 11
0 33 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 66 239 0 10 11
0 31 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 67 151 0 10 11
0 34 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 69 96 0 1 11
0 32
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 70 45 0 1 11
0 30
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 793 607 0 3 22
0 4 5 3
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6B
-13 -4 8 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
8901 0 0
2
43337.5 0
0
9 2-In XOR~
219 786 558 0 3 22
0 4 5 2
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U8A
0 -3 21 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
7361 0 0
2
43337.5 0
0
9 2-In AND~
219 795 508 0 3 22
0 8 7 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6A
-13 -3 8 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
4747 0 0
2
43337.5 0
0
9 2-In XOR~
219 788 460 0 3 22
0 7 8 5
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U5D
0 -3 21 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
972 0 0
2
43337.5 0
0
9 2-In AND~
219 572 706 0 3 22
0 9 10 4
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4D
-13 -3 8 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
3472 0 0
2
43337.5 0
0
9 2-In XOR~
219 565 659 0 3 22
0 10 9 11
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U5C
-1 -3 20 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
9998 0 0
2
43337.5 0
0
9 2-In AND~
219 572 607 0 3 22
0 14 13 12
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4C
-13 -4 8 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
3536 0 0
2
43337.5 0
0
9 2-In XOR~
219 565 558 0 3 22
0 14 13 9
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U5B
-1 -4 20 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
4597 0 0
2
43337.5 0
0
9 2-In AND~
219 574 514 0 3 22
0 16 17 15
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-13 -3 8 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
3835 0 0
2
43337.5 0
0
9 2-In XOR~
219 568 465 0 3 22
0 16 17 13
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U5A
0 -4 21 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
3670 0 0
2
43337.5 0
0
9 2-In AND~
219 357 707 0 3 22
0 19 20 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-13 -4 8 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
5616 0 0
2
43337.5 0
0
9 2-In XOR~
219 351 659 0 3 22
0 19 20 18
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U2D
1 -3 22 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
9323 0 0
2
43337.5 0
0
9 2-In AND~
219 359 605 0 3 22
0 22 23 21
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U11D
-16 -3 12 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
317 0 0
2
43337.5 0
0
9 2-In XOR~
219 353 559 0 3 22
0 22 23 19
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U2C
0 -4 21 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
3108 0 0
2
43337.5 0
0
9 2-In AND~
219 361 513 0 3 22
0 25 26 24
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U11C
-16 -4 12 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
4299 0 0
2
43337.5 0
0
9 2-In XOR~
219 355 469 0 3 22
0 25 26 22
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U2B
0 -4 21 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
9672 0 0
2
43337.5 0
0
9 2-In AND~
219 197 515 0 3 22
0 27 28 23
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U11B
-15 -4 13 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
7876 0 0
2
43337.5 0
0
9 2-In XOR~
219 190 471 0 3 22
0 27 28 36
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U2A
0 -4 21 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
6369 0 0
2
43337.5 0
0
14 Logic Display~
6 963 755 0 1 2
10 29
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9172 0 0
2
5.89859e-315 0
0
14 Logic Display~
6 851 755 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7100 0 0
2
5.89859e-315 0
0
14 Logic Display~
6 643 755 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3820 0 0
2
5.89859e-315 0
0
14 Logic Display~
6 433 755 0 1 2
10 18
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7678 0 0
2
5.89859e-315 0
0
14 Logic Display~
6 260 754 0 1 2
10 36
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
961 0 0
2
5.89859e-315 0
0
14 Logic Display~
6 145 755 0 1 2
10 37
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3178 0 0
2
5.89859e-315 0
0
8 2-In OR~
219 873 506 0 3 22
0 6 3 29
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7C
-1 -4 20 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
3409 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 789 394 0 3 22
0 30 31 8
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U11A
-15 -11 13 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3951 0 0
2
5.89859e-315 0
0
8 2-In OR~
219 665 511 0 3 22
0 15 12 7
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7B
-1 -4 20 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
8885 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 587 394 0 3 22
0 31 32 10
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3D
-12 -11 9 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
3780 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 549 395 0 3 22
0 33 30 14
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3C
-12 -11 9 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
9265 0 0
2
5.89859e-315 0
0
8 2-In OR~
219 441 513 0 3 22
0 24 21 17
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7A
-1 -4 20 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
9442 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 398 396 0 3 22
0 31 34 20
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3B
-12 -11 9 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
9424 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 358 396 0 3 22
0 33 32 26
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3A
-12 -11 9 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
9968 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 317 397 0 3 22
0 35 30 25
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1D
-12 -11 9 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
9281 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 213 396 0 3 22
0 33 34 28
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1C
-12 -11 9 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
8464 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 169 396 0 3 22
0 35 32 27
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1B
-12 -10 9 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
7168 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 121 397 0 3 22
0 34 35 37
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1A
-12 -10 9 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3171 0 0
2
5.89859e-315 0
0
72
3 1 2 0 0 8320 0 8 26 0 0 5
819 558
834 558
834 782
851 782
851 773
3 2 3 0 0 8320 0 7 31 0 0 4
814 607
845 607
845 515
860 515
0 1 4 0 0 8192 0 0 7 5 0 3
713 549
713 598
769 598
0 2 5 0 0 4096 0 0 7 6 0 3
738 567
738 616
769 616
3 1 4 0 0 8320 0 11 8 0 0 4
593 706
655 706
655 549
770 549
3 2 5 0 0 12416 0 10 8 0 0 6
821 460
833 460
833 533
738 533
738 567
770 567
3 1 6 0 0 12416 0 9 31 0 0 4
816 508
827 508
827 497
860 497
0 2 7 0 0 4096 0 0 9 11 0 3
727 451
727 517
771 517
0 1 8 0 0 8192 0 0 9 10 0 3
714 469
714 499
771 499
3 2 8 0 0 8320 0 32 10 0 0 5
787 417
787 430
714 430
714 469
772 469
3 1 7 0 0 8320 0 33 10 0 0 3
698 511
698 451
772 451
0 1 9 0 0 4096 0 0 11 16 0 3
524 667
524 697
548 697
0 2 10 0 0 4096 0 0 11 15 0 3
517 648
517 715
548 715
3 1 11 0 0 8320 0 12 27 0 0 5
598 659
626 659
626 782
643 782
643 773
3 1 10 0 0 12416 0 34 12 0 0 7
585 417
585 426
603 426
603 639
517 639
517 650
549 650
3 2 9 0 0 12416 0 14 12 0 0 6
598 558
618 558
618 632
524 632
524 668
549 668
3 2 12 0 0 8320 0 13 33 0 0 4
593 607
626 607
626 520
652 520
0 2 13 0 0 4096 0 0 13 21 0 3
517 567
517 616
548 616
0 1 14 0 0 4096 0 0 13 20 0 3
510 549
510 598
548 598
3 1 14 0 0 8320 0 35 14 0 0 4
547 418
510 418
510 549
549 549
3 2 13 0 0 12416 0 16 14 0 0 6
601 465
611 465
611 536
517 536
517 567
549 567
3 1 15 0 0 4224 0 15 33 0 0 4
595 514
626 514
626 502
652 502
0 1 16 0 0 4096 0 0 15 25 0 3
530 456
530 505
550 505
0 2 17 0 0 4224 0 0 15 26 0 3
517 474
517 523
550 523
3 1 16 0 0 8320 0 17 16 0 0 4
378 707
494 707
494 456
552 456
3 2 17 0 0 0 0 36 16 0 0 4
474 513
503 513
503 474
552 474
3 1 18 0 0 8320 0 18 28 0 0 5
384 659
412 659
412 782
433 782
433 773
0 1 19 0 0 8192 0 0 17 30 0 3
283 654
283 698
333 698
0 2 20 0 0 4096 0 0 17 31 0 3
292 672
292 716
333 716
3 1 19 0 0 12416 0 20 18 0 0 8
386 559
404 559
404 628
283 628
283 654
283 654
283 650
335 650
3 2 20 0 0 4224 0 37 18 0 0 7
396 419
396 635
292 635
292 672
292 672
292 668
335 668
3 2 21 0 0 8320 0 19 36 0 0 4
380 605
412 605
412 522
428 522
0 1 22 0 0 4096 0 0 19 36 0 3
300 549
300 596
335 596
0 2 23 0 0 4096 0 0 19 35 0 3
292 568
292 614
335 614
3 2 23 0 0 4224 0 23 20 0 0 4
218 515
292 515
292 568
337 568
3 1 22 0 0 12416 0 22 20 0 0 6
388 469
404 469
404 536
300 536
300 550
337 550
3 1 24 0 0 4224 0 21 36 0 0 4
382 513
412 513
412 504
428 504
0 1 25 0 0 4224 0 0 21 40 0 3
315 460
315 504
337 504
0 2 26 0 0 4096 0 0 21 41 0 3
300 478
300 522
337 522
3 1 25 0 0 0 0 39 22 0 0 3
315 420
315 460
339 460
3 2 26 0 0 8320 0 38 22 0 0 5
356 419
356 439
300 439
300 478
339 478
0 1 27 0 0 4224 0 0 23 44 0 3
167 461
167 506
173 506
0 2 28 0 0 4096 0 0 23 45 0 3
152 480
152 524
173 524
3 1 27 0 0 0 0 41 24 0 0 3
167 419
167 462
174 462
3 2 28 0 0 8320 0 40 24 0 0 5
211 419
211 440
152 440
152 480
174 480
3 1 29 0 0 8320 0 31 25 0 0 7
906 506
947 506
947 774
951 774
951 781
963 781
963 773
1 0 30 0 0 4096 0 32 0 0 72 2
796 372
796 45
2 0 31 0 0 4096 0 32 0 0 69 2
778 372
778 239
1 0 31 0 0 0 0 34 0 0 69 2
594 372
594 239
2 0 32 0 0 4096 0 34 0 0 71 2
576 372
576 96
1 0 33 0 0 4096 0 35 0 0 68 2
556 373
556 294
2 0 30 0 0 4096 0 35 0 0 72 2
538 373
538 45
1 0 31 0 0 4096 0 37 0 0 69 2
405 374
405 239
2 0 34 0 0 4096 0 37 0 0 70 2
387 374
387 151
1 0 33 0 0 4096 0 38 0 0 68 2
365 374
365 294
2 0 32 0 0 4096 0 38 0 0 71 2
347 374
347 96
1 0 35 0 0 4096 0 39 0 0 67 2
324 375
324 353
2 0 30 0 0 4096 0 39 0 0 72 2
306 375
306 45
3 1 36 0 0 8320 0 24 29 0 0 7
223 471
236 471
236 773
248 773
248 780
260 780
260 772
1 0 33 0 0 0 0 40 0 0 68 2
220 374
220 294
2 0 34 0 0 0 0 40 0 0 70 2
202 374
202 151
1 0 35 0 0 0 0 41 0 0 67 2
176 374
176 353
2 0 32 0 0 0 0 41 0 0 71 2
158 374
158 96
3 1 37 0 0 4224 0 42 30 0 0 6
119 420
119 773
133 773
133 781
145 781
145 773
1 0 34 0 0 4096 0 42 0 0 70 2
128 375
128 151
2 0 35 0 0 0 0 42 0 0 67 2
110 375
110 353
1 0 35 0 0 4224 0 1 0 0 0 2
75 353
1156 353
1 0 33 0 0 4224 0 2 0 0 0 2
76 294
1155 294
1 0 31 0 0 4224 0 3 0 0 0 2
78 239
1156 239
1 0 34 0 0 4224 0 4 0 0 0 2
79 151
1156 151
1 0 32 0 0 4224 0 5 0 0 0 2
81 96
1155 96
1 0 30 0 0 4224 0 6 0 0 0 2
82 45
1155 45
12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
20 23 57 47
30 31 46 47
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
20 74 57 98
30 82 46 98
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
19 127 56 151
29 135 45 151
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
18 215 55 239
28 223 44 239
2 B2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
17 273 54 297
27 281 43 297
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
16 329 53 353
26 337 42 353
2 B0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
127 702 164 726
137 710 153 726
2 SO
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
242 702 279 726
252 710 268 726
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
415 703 452 727
425 711 441 727
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
624 705 661 729
634 713 650 729
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
833 704 870 728
843 712 859 728
2 S4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
944 702 981 726
954 710 970 726
2 S5
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
