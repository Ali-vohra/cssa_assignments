CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 80 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
16
13 Logic Switch~
5 113 340 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
969 0 0
2
5.89865e-315 0
0
13 Logic Switch~
5 114 295 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8402 0 0
2
5.89865e-315 0
0
13 Logic Switch~
5 113 183 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3751 0 0
2
5.89865e-315 0
0
13 Logic Switch~
5 113 131 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4292 0 0
2
5.89865e-315 0
0
14 Logic Display~
6 799 774 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6118 0 0
2
5.89865e-315 0
0
14 Logic Display~
6 650 775 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
34 0 0
2
5.89865e-315 0
0
7 Ground~
168 824 151 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6357 0 0
2
5.89865e-315 0
0
7 Ground~
168 664 153 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
319 0 0
2
5.89865e-315 0
0
6 Diode~
219 709 413 0 2 5
0 5 6
0
0 0 848 0
6 1N1185
-21 -18 21 -10
2 D6
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
9 DOIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
3976 0 0
2
5.89865e-315 0
0
6 Diode~
219 565 416 0 2 5
0 5 3
0
0 0 848 0
6 1N1185
-21 -18 21 -10
2 D5
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
9 DOIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
7634 0 0
2
5.89865e-315 0
0
6 Diode~
219 565 510 0 2 5
0 4 3
0
0 0 848 0
6 1N1185
-21 -18 21 -10
2 D3
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
9 DOIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
523 0 0
2
5.89865e-315 0
0
6 Diode~
219 564 324 0 2 5
0 7 3
0
0 0 848 0
6 1N1185
-21 -18 21 -10
2 D2
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
9 DOIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
6748 0 0
2
5.89865e-315 0
0
6 Diode~
219 710 240 0 2 5
0 8 6
0
0 0 848 0
6 1N1185
-21 -18 21 -10
2 D1
-7 -28 7 -20
0
0
11 %D %1 %2 %M
0
0
9 DOIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
6901 0 0
2
5.89865e-315 0
0
8 2-4 DEC~
94 328 292 0 8 17
0 12 11 10 9 4 5 7 8
8 2-4 DEC~
1 0 560 0
7 2-4 DEC
-21 -77 28 -69
2 U1
-3 -77 11 -69
0
0
0
0
0
0
17

0 1 2 7 8 11 12 13 14 1
2 7 8 11 12 13 14 0
0 0 0 0 1 0 0 0
1 U
842 0 0
2
5.89861e-315 0
0
9 Resistor~
219 607 155 0 4 5
0 3 2 0 -1
0
0 0 880 90
2 1k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3277 0 0
2
5.89865e-315 0
0
9 Resistor~
219 753 157 0 4 5
0 6 2 0 -1
0
0 0 880 90
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4212 0 0
2
5.89865e-315 0
0
22
2 0 3 0 0 4096 0 11 0 0 12 2
575 510
607 510
1 0 4 0 0 8192 0 11 0 0 3 3
555 510
523 510
523 546
5 0 4 0 0 12416 0 14 0 0 0 4
378 319
420 319
420 546
1135 546
2 0 3 0 0 0 0 10 0 0 12 2
575 416
607 416
1 0 5 0 0 8192 0 9 0 0 8 3
699 413
671 413
671 455
2 0 6 0 0 4096 0 9 0 0 11 2
719 413
753 413
1 0 5 0 0 0 0 10 0 0 8 3
555 416
523 416
523 455
6 0 5 0 0 12416 0 14 0 0 0 4
378 305
411 305
411 455
1135 455
2 0 3 0 0 4096 0 12 0 0 12 2
574 324
607 324
2 0 6 0 0 0 0 13 0 0 11 2
720 240
753 240
1 1 6 0 0 4224 0 16 5 0 0 6
753 175
753 502
752 502
752 797
799 797
799 792
1 1 3 0 0 4224 0 15 6 0 0 4
607 173
607 797
650 797
650 793
1 0 7 0 0 8192 0 12 0 0 14 3
554 324
524 324
524 363
7 0 7 0 0 12416 0 14 0 0 0 4
378 292
402 292
402 363
1135 363
2 1 2 0 0 8320 0 16 7 0 0 4
753 139
753 135
824 135
824 145
2 1 2 0 0 0 0 15 8 0 0 4
607 137
607 133
664 133
664 147
1 0 8 0 0 8192 0 13 0 0 18 3
700 240
676 240
676 279
8 0 8 0 0 4224 0 14 0 0 0 2
378 279
1134 279
1 4 9 0 0 8320 0 1 14 0 0 3
125 340
125 346
286 346
1 3 10 0 0 4224 0 2 14 0 0 4
126 295
234 295
234 332
286 332
1 2 11 0 0 4224 0 3 14 0 0 4
125 183
234 183
234 265
286 265
1 1 12 0 0 8320 0 4 14 0 0 4
125 131
223 131
223 252
286 252
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
55 112 92 136
65 120 81 136
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
54 162 91 186
64 170 80 186
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
57 279 94 303
67 287 83 303
2 E2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
55 317 92 341
65 325 81 341
2 E1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
631 700 668 724
641 708 657 724
2 F1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
780 701 817 725
790 709 806 725
2 F2
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
