CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
60 10 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
30
13 Logic Switch~
5 79 484 0 1 11
0 6
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 77 420 0 1 11
0 5
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 78 350 0 1 11
0 14
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 76 201 0 1 11
0 18
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 72 140 0 1 11
0 20
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 72 73 0 1 11
0 27
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
5.89855e-315 0
0
9 Inverter~
13 126 469 0 2 22
0 6 13
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 4 0
1 U
8901 0 0
2
5.89855e-315 0
0
9 Inverter~
13 124 402 0 2 22
0 5 12
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 4 0
1 U
7361 0 0
2
5.89855e-315 0
0
9 Inverter~
13 123 331 0 2 22
0 14 7
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 4 0
1 U
4747 0 0
2
5.89855e-315 0
0
5 4073~
219 423 481 0 4 22
0 4 3 2 28
0
0 0 608 0
4 4073
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 512 3 2 2 0
1 U
972 0 0
2
5.89855e-315 0
0
5 4082~
219 426 371 0 5 22
0 11 10 9 8 29
0
0 0 608 0
4 4082
-7 -24 21 -16
3 U9A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 512 2 1 9 0
1 U
3472 0 0
2
5.89855e-315 0
0
5 4071~
219 289 517 0 3 22
0 6 5 2
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U8C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 8 0
1 U
9998 0 0
2
5.89855e-315 0
0
5 4071~
219 289 451 0 3 22
0 7 5 4
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U8B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 8 0
1 U
3536 0 0
2
5.89855e-315 0
0
5 4071~
219 292 377 0 3 22
0 7 6 3
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U8A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 8 0
1 U
4597 0 0
2
5.89855e-315 0
0
8 3-In OR~
219 184 538 0 4 22
0 6 7 12 8
0
0 0 608 0
4 4075
-14 -24 14 -16
3 U7B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 7 0
1 U
3835 0 0
2
5.89855e-315 0
0
8 3-In OR~
219 185 476 0 4 22
0 7 5 13 9
0
0 0 608 0
4 4075
-14 -24 14 -16
3 U7A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 7 0
1 U
3670 0 0
2
5.89855e-315 0
0
8 3-In OR~
219 187 415 0 4 22
0 14 12 13 10
0
0 0 608 0
4 4075
-14 -24 14 -16
3 U6C
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 6 0
1 U
5616 0 0
2
5.89855e-315 0
0
8 3-In OR~
219 188 351 0 4 22
0 14 5 6 11
0
0 0 608 0
4 4075
-14 -24 14 -16
3 U6B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 6 0
1 U
9323 0 0
2
5.89855e-315 0
0
8 3-In OR~
219 424 170 0 4 22
0 15 16 17 30
0
0 0 608 0
4 4075
-14 -24 14 -16
3 U6A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 512 3 1 6 0
1 U
317 0 0
2
5.89855e-315 0
0
8 4-In OR~
219 426 81 0 5 22
0 24 23 22 21 31
0
0 0 608 0
4 4072
-14 -24 14 -16
3 U5A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 512 2 1 5 0
1 U
3108 0 0
2
5.89855e-315 0
0
9 Inverter~
13 116 186 0 2 22
0 18 25
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 4 0
1 U
4299 0 0
2
5.89855e-315 0
0
9 Inverter~
13 116 123 0 2 22
0 20 26
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
9672 0 0
2
5.89855e-315 0
0
9 Inverter~
13 116 56 0 2 22
0 27 19
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
7876 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 310 203 0 3 22
0 19 18 17
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
6369 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 313 138 0 3 22
0 20 18 16
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
9172 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 312 67 0 3 22
0 19 20 15
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
7100 0 0
2
5.89855e-315 0
0
5 4073~
219 198 234 0 4 22
0 27 26 25 21
0
0 0 608 0
4 4073
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 2 0
1 U
3820 0 0
2
5.89855e-315 0
0
5 4073~
219 199 171 0 4 22
0 19 20 25 22
0
0 0 608 0
4 4073
-7 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 1 0
1 U
7678 0 0
2
5.89855e-315 0
0
5 4073~
219 201 108 0 4 22
0 19 26 18 23
0
0 0 608 0
4 4073
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 1 0
1 U
961 0 0
2
5.89855e-315 0
0
5 4073~
219 201 44 0 4 22
0 27 20 18 24
0
0 0 608 0
4 4073
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 1 0
1 U
3178 0 0
2
5.89855e-315 0
0
56
3 3 2 0 0 4224 0 12 10 0 0 4
322 517
391 517
391 490
399 490
3 2 3 0 0 8320 0 14 10 0 0 4
325 377
376 377
376 481
399 481
3 1 4 0 0 4224 0 13 10 0 0 4
322 451
381 451
381 472
399 472
1 2 5 0 0 8320 0 2 12 0 0 6
89 420
152 420
152 558
268 558
268 526
276 526
1 1 6 0 0 12288 0 1 12 0 0 4
91 484
168 484
168 508
276 508
1 2 5 0 0 0 0 2 13 0 0 6
89 420
153 420
153 496
268 496
268 460
276 460
2 1 7 0 0 4096 0 9 13 0 0 4
144 331
268 331
268 442
276 442
1 2 6 0 0 12416 0 1 14 0 0 4
91 484
153 484
153 386
279 386
2 1 7 0 0 4096 0 9 14 0 0 4
144 331
271 331
271 368
279 368
4 4 8 0 0 4224 0 15 11 0 0 4
217 538
384 538
384 385
402 385
4 3 9 0 0 4224 0 16 11 0 0 4
218 476
389 476
389 376
402 376
4 2 10 0 0 4224 0 17 11 0 0 4
220 415
394 415
394 367
402 367
4 1 11 0 0 4224 0 18 11 0 0 4
221 351
394 351
394 358
402 358
2 3 12 0 0 8320 0 8 15 0 0 4
145 402
153 402
153 547
171 547
2 2 7 0 0 8320 0 9 15 0 0 4
144 331
153 331
153 538
172 538
1 1 6 0 0 0 0 1 15 0 0 4
91 484
153 484
153 529
171 529
2 3 13 0 0 8192 0 7 16 0 0 4
147 469
159 469
159 485
172 485
1 2 5 0 0 0 0 2 16 0 0 4
89 420
154 420
154 476
173 476
2 1 7 0 0 0 0 9 16 0 0 4
144 331
159 331
159 467
172 467
2 3 13 0 0 8320 0 7 17 0 0 4
147 469
166 469
166 424
174 424
2 2 12 0 0 0 0 8 17 0 0 4
145 402
151 402
151 415
175 415
1 1 14 0 0 4096 0 3 17 0 0 4
90 350
156 350
156 406
174 406
1 1 6 0 0 0 0 1 7 0 0 4
91 484
103 484
103 469
111 469
1 1 5 0 0 0 0 2 8 0 0 4
89 420
101 420
101 402
109 402
1 1 14 0 0 0 0 3 9 0 0 4
90 350
100 350
100 331
108 331
1 3 6 0 0 0 0 1 18 0 0 4
91 484
162 484
162 360
175 360
1 2 5 0 0 0 0 2 18 0 0 4
89 420
167 420
167 351
176 351
1 1 14 0 0 4224 0 3 18 0 0 4
90 350
167 350
167 342
175 342
3 1 15 0 0 8320 0 26 19 0 0 4
333 67
388 67
388 161
411 161
3 2 16 0 0 4224 0 25 19 0 0 4
334 138
403 138
403 170
412 170
3 3 17 0 0 4224 0 24 19 0 0 4
331 203
403 203
403 179
411 179
1 2 18 0 0 4096 0 4 24 0 0 4
88 201
278 201
278 212
286 212
2 1 19 0 0 12416 0 23 24 0 0 4
137 56
145 56
145 194
286 194
1 2 18 0 0 4224 0 4 25 0 0 4
88 201
281 201
281 147
289 147
1 1 20 0 0 4096 0 5 25 0 0 4
84 140
276 140
276 129
289 129
1 2 20 0 0 4224 0 5 26 0 0 4
84 140
280 140
280 76
288 76
2 1 19 0 0 0 0 23 26 0 0 6
137 56
173 56
173 64
280 64
280 58
288 58
4 4 21 0 0 4224 0 27 20 0 0 4
219 234
391 234
391 95
409 95
4 3 22 0 0 4224 0 28 20 0 0 4
220 171
396 171
396 86
409 86
4 2 23 0 0 4224 0 29 20 0 0 4
222 108
401 108
401 77
409 77
4 1 24 0 0 4224 0 30 20 0 0 4
222 44
401 44
401 68
409 68
2 3 25 0 0 8320 0 21 27 0 0 4
137 186
146 186
146 243
174 243
2 2 26 0 0 8320 0 22 27 0 0 4
137 123
141 123
141 234
174 234
1 1 27 0 0 8320 0 6 27 0 0 4
84 73
151 73
151 225
174 225
2 3 25 0 0 0 0 21 28 0 0 4
137 186
167 186
167 180
175 180
1 2 20 0 0 0 0 5 28 0 0 4
84 140
167 140
167 171
175 171
2 1 19 0 0 0 0 23 28 0 0 4
137 56
147 56
147 162
175 162
1 3 18 0 0 0 0 4 29 0 0 4
88 201
154 201
154 117
177 117
2 2 26 0 0 0 0 22 29 0 0 4
137 123
169 123
169 108
177 108
2 1 19 0 0 0 0 23 29 0 0 4
137 56
154 56
154 99
177 99
1 1 18 0 0 0 0 4 21 0 0 4
88 201
93 201
93 186
101 186
1 1 20 0 0 0 0 5 22 0 0 4
84 140
93 140
93 123
101 123
1 1 27 0 0 0 0 6 23 0 0 4
84 73
93 73
93 56
101 56
1 3 18 0 0 0 0 4 30 0 0 4
88 201
159 201
159 53
177 53
1 2 20 0 0 0 0 5 30 0 0 4
84 140
164 140
164 44
177 44
1 1 27 0 0 0 0 6 30 0 0 4
84 73
169 73
169 35
177 35
7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
157 579 298 603
167 587 287 603
15 FULL SUBTRACTOR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
454 64 555 88
464 72 544 88
10 Difference
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
450 157 519 181
460 165 508 181
6 Borrow
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
442 355 543 379
452 363 532 379
10 Difference
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
437 467 506 491
447 475 495 491
6 Borrow
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
547 111 632 135
557 119 621 135
8 SOP Form
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
564 413 649 437
574 421 638 437
8 POS Form
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
