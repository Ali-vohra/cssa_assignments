CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
30 40 30 130 10
176 80 1534 843
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
31
13 Logic Switch~
5 92 430 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89857e-315 0
0
13 Logic Switch~
5 94 391 0 1 11
0 21
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.89857e-315 0
0
13 Logic Switch~
5 94 300 0 1 11
0 22
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3124 0 0
2
5.89857e-315 0
0
13 Logic Switch~
5 95 259 0 1 11
0 25
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
5.89857e-315 0
0
13 Logic Switch~
5 93 165 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.89857e-315 0
0
13 Logic Switch~
5 92 123 0 10 11
0 29 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
5.89857e-315 0
0
14 Logic Display~
6 934 357 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8901 0 0
2
5.89857e-315 0
0
14 Logic Display~
6 930 222 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7361 0 0
2
5.89857e-315 0
0
14 Logic Display~
6 930 70 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4747 0 0
2
5.89857e-315 0
0
5 4073~
219 710 254 0 4 22
0 7 6 5 3
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 5 0
1 U
972 0 0
2
5.89857e-315 0
0
8 3-In OR~
219 710 387 0 4 22
0 10 9 8 2
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U6B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 6 0
1 U
3472 0 0
2
5.89857e-315 0
0
8 3-In OR~
219 705 115 0 4 22
0 15 14 13 4
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U6A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 6 0
1 U
9998 0 0
2
5.89857e-315 0
0
9 2-In AND~
219 526 359 0 3 22
0 7 12 10
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
3536 0 0
2
5.89857e-315 0
0
5 4073~
219 525 420 0 4 22
0 7 6 11 9
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 5 0
1 U
4597 0 0
2
5.89857e-315 0
0
5 4073~
219 527 156 0 4 22
0 7 6 16 13
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 5 0
1 U
3835 0 0
2
5.89857e-315 0
0
9 2-In AND~
219 526 101 0 3 22
0 7 17 14
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
3670 0 0
2
5.89857e-315 0
0
9 2-In AND~
219 378 426 0 3 22
0 19 18 11
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
5616 0 0
2
5.89857e-315 0
0
9 2-In AND~
219 378 378 0 3 22
0 21 20 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
9323 0 0
2
5.89857e-315 0
0
9 2-In AND~
219 377 298 0 3 22
0 23 22 12
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
317 0 0
2
5.89857e-315 0
0
9 2-In AND~
219 378 244 0 3 22
0 25 24 17
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
3108 0 0
2
5.89857e-315 0
0
9 2-In AND~
219 377 151 0 3 22
0 27 26 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
4299 0 0
2
5.89857e-315 0
0
9 2-In AND~
219 375 102 0 3 22
0 29 28 15
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
9672 0 0
2
5.89857e-315 0
0
9 Inverter~
13 186 427 0 2 22
0 18 20
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
7876 0 0
2
5.89857e-315 0
0
9 Inverter~
13 185 386 0 2 22
0 21 19
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 2 0
1 U
6369 0 0
2
5.89857e-315 0
0
9 Inverter~
13 184 291 0 2 22
0 22 24
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
9172 0 0
2
5.89857e-315 0
0
9 Inverter~
13 182 255 0 2 22
0 25 23
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
7100 0 0
2
5.89857e-315 0
0
9 Inverter~
13 178 151 0 2 22
0 26 28
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
3820 0 0
2
5.89857e-315 0
0
9 Inverter~
13 177 116 0 2 22
0 29 27
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
7678 0 0
2
5.89857e-315 0
0
10 2-In XNOR~
219 260 398 0 3 22
0 21 18 5
0
0 0 624 0
4 4077
-7 -24 21 -16
3 U1C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 1 0
1 U
961 0 0
2
5.89857e-315 0
0
10 2-In XNOR~
219 265 270 0 3 22
0 25 22 6
0
0 0 624 0
4 4077
-7 -24 21 -16
3 U1B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
3178 0 0
2
5.89857e-315 0
0
10 2-In XNOR~
219 266 124 0 3 22
0 29 26 7
0
0 0 624 0
4 4077
-7 -24 21 -16
3 U1A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
3409 0 0
2
5.89857e-315 0
0
46
4 1 2 0 0 4224 0 11 7 0 0 3
743 387
934 387
934 375
4 1 3 0 0 4224 0 10 8 0 0 3
731 254
930 254
930 240
4 1 4 0 0 4224 0 12 9 0 0 3
738 115
930 115
930 88
3 3 5 0 0 4224 0 29 10 0 0 4
299 398
673 398
673 263
686 263
3 2 6 0 0 4224 0 30 10 0 0 4
304 270
678 270
678 254
686 254
3 1 7 0 0 4224 0 31 10 0 0 4
305 124
678 124
678 245
686 245
3 3 8 0 0 8320 0 21 11 0 0 4
398 151
482 151
482 396
697 396
4 2 9 0 0 4224 0 14 11 0 0 4
546 420
689 420
689 387
698 387
3 1 10 0 0 4224 0 13 11 0 0 4
547 359
689 359
689 378
697 378
3 3 11 0 0 4224 0 17 14 0 0 4
399 426
493 426
493 429
501 429
3 2 6 0 0 0 0 30 14 0 0 4
304 270
488 270
488 420
501 420
3 1 7 0 0 0 0 31 14 0 0 4
305 124
473 124
473 411
501 411
3 2 12 0 0 4224 0 19 13 0 0 4
398 298
494 298
494 368
502 368
3 1 7 0 0 0 0 31 13 0 0 4
305 124
479 124
479 350
502 350
4 3 13 0 0 4224 0 15 12 0 0 4
548 156
684 156
684 124
692 124
3 2 14 0 0 4224 0 16 12 0 0 4
547 101
679 101
679 115
693 115
3 1 15 0 0 12416 0 22 12 0 0 6
396 102
498 102
498 121
684 121
684 106
692 106
3 3 16 0 0 8320 0 18 15 0 0 4
399 378
485 378
485 165
503 165
3 2 6 0 0 0 0 30 15 0 0 4
304 270
495 270
495 156
503 156
3 1 7 0 0 0 0 31 15 0 0 4
305 124
485 124
485 147
503 147
3 2 17 0 0 8320 0 20 16 0 0 4
399 244
489 244
489 110
502 110
3 1 7 0 0 0 0 31 16 0 0 4
305 124
494 124
494 92
502 92
1 2 18 0 0 12416 0 1 17 0 0 6
104 430
157 430
157 442
346 442
346 435
354 435
2 1 19 0 0 12416 0 24 17 0 0 4
206 386
240 386
240 417
354 417
2 2 20 0 0 4224 0 23 18 0 0 4
207 427
346 427
346 387
354 387
1 1 21 0 0 12416 0 2 18 0 0 4
106 391
156 391
156 369
354 369
1 2 22 0 0 12416 0 3 19 0 0 4
106 300
155 300
155 307
353 307
2 1 23 0 0 12416 0 26 19 0 0 4
203 255
245 255
245 289
353 289
2 2 24 0 0 4224 0 25 20 0 0 4
205 291
346 291
346 253
354 253
1 1 25 0 0 12416 0 4 20 0 0 4
107 259
153 259
153 235
354 235
1 2 26 0 0 4224 0 5 21 0 0 4
105 165
345 165
345 160
353 160
2 1 27 0 0 12416 0 28 21 0 0 4
198 116
246 116
246 142
353 142
2 2 28 0 0 4224 0 27 22 0 0 4
199 151
343 151
343 111
351 111
1 1 29 0 0 12416 0 6 22 0 0 4
104 123
148 123
148 93
351 93
1 1 18 0 0 0 0 1 23 0 0 4
104 430
163 430
163 427
171 427
1 1 21 0 0 0 0 2 24 0 0 4
106 391
162 391
162 386
170 386
1 1 22 0 0 0 0 3 25 0 0 4
106 300
161 300
161 291
169 291
1 1 25 0 0 0 0 4 26 0 0 4
107 259
159 259
159 255
167 255
1 1 26 0 0 0 0 5 27 0 0 4
105 165
155 165
155 151
163 151
1 1 29 0 0 0 0 6 28 0 0 5
104 123
104 117
154 117
154 116
162 116
1 2 18 0 0 0 0 1 29 0 0 4
104 430
167 430
167 407
244 407
1 1 21 0 0 0 0 2 29 0 0 6
106 391
166 391
166 401
236 401
236 389
244 389
1 2 22 0 0 0 0 3 30 0 0 6
106 300
165 300
165 276
241 276
241 279
249 279
1 1 25 0 0 0 0 4 30 0 0 6
107 259
163 259
163 270
241 270
241 261
249 261
1 2 26 0 0 0 0 5 31 0 0 4
105 165
242 165
242 133
250 133
1 1 29 0 0 0 0 6 31 0 0 6
104 123
158 123
158 101
242 101
242 115
250 115
10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
39 103 76 127
49 111 65 127
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
37 140 74 164
47 148 63 164
2 B2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
35 235 72 259
45 243 61 259
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
34 283 71 307
44 291 60 307
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
37 370 74 394
47 378 63 394
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
36 414 73 438
46 422 62 438
2 B0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
946 62 991 86
956 70 980 86
3 A>B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
948 208 993 232
958 216 982 232
3 A=B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
949 345 994 369
959 353 983 369
3 A<B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
495 488 644 512
505 496 633 512
16 3 BIT COMPARATOR
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
