CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 110 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
27
13 Logic Switch~
5 472 315 0 10 11
0 29 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43331 0
0
9 2-In AND~
219 695 212 0 3 22
0 4 3 2
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
391 0 0
2
43331.1 0
0
9 Inverter~
13 702 290 0 2 22
0 5 4
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U7A
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 5 0
1 U
3124 0 0
2
43331.1 0
0
9 Inverter~
13 705 416 0 2 22
0 6 3
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U4F
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
3421 0 0
2
43331.1 0
0
5 4073~
219 625 308 0 4 22
0 9 7 8 5
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 4 0
1 U
8157 0 0
2
43331.1 0
0
9 Inverter~
13 568 393 0 2 22
0 10 8
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 2 0
1 U
5572 0 0
2
43331.1 0
0
9 Inverter~
13 570 234 0 2 22
0 11 9
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
8901 0 0
2
43331.1 0
0
8 4-In OR~
219 522 393 0 5 22
0 15 14 13 12 10
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U5B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 3 0
1 U
7361 0 0
2
43331.1 0
0
8 4-In OR~
219 523 234 0 5 22
0 19 18 17 16 11
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U5A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 3 0
1 U
4747 0 0
2
43331.1 0
0
9 Inverter~
13 600 434 0 2 22
0 7 6
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
972 0 0
2
43331.1 0
0
14 Logic Display~
6 804 211 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3472 0 0
2
43331.1 0
0
14 Logic Display~
6 804 312 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9998 0 0
2
43331.1 0
0
14 Logic Display~
6 805 403 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3536 0 0
2
43331.1 0
0
9 Inverter~
13 339 501 0 2 22
0 45 38
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
4597 0 0
2
43331 0
0
9 Inverter~
13 339 464 0 2 22
0 44 39
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
3835 0 0
2
43331 0
0
9 Inverter~
13 339 428 0 2 22
0 43 40
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
3670 0 0
2
43331 0
0
9 Inverter~
13 339 396 0 2 22
0 42 41
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
5616 0 0
2
43331 0
0
9 Inverter~
13 339 330 0 2 22
0 34 30
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
9323 0 0
2
43331 0
0
9 Inverter~
13 339 297 0 2 22
0 35 31
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
317 0 0
2
43331 0
0
9 Inverter~
13 338 264 0 2 22
0 36 32
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
3108 0 0
2
43331 0
0
9 Inverter~
13 338 231 0 2 22
0 37 33
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
4299 0 0
2
43331 0
0
6 74LS83
105 475 389 0 14 29
0 20 21 22 23 41 40 39 38 24
15 14 13 12 7
0
0 0 4848 0
5 74F83
-18 -60 17 -52
2 U2
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 0 0 0 0
1 U
9672 0 0
2
43331 0
0
6 74LS83
105 476 230 0 14 29
0 25 26 27 28 33 32 31 30 29
19 18 17 16 24
0
0 0 4848 0
5 74F83
-18 -60 17 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 0 0 0 0
1 U
7876 0 0
2
43331 0
0
8 Hex Key~
166 256 86 0 11 12
0 34 35 36 37 0 0 0 0 0
13 68
0
0 0 4656 0
0
4 KPD4
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
6369 0 0
2
43331 0
0
8 Hex Key~
166 213 86 0 11 12
0 45 44 43 42 0 0 0 0 0
3 51
0
0 0 4656 0
0
4 KPD3
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
9172 0 0
2
43331 0
0
8 Hex Key~
166 97 87 0 11 12
0 28 27 26 25 0 0 0 0 0
13 68
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
7100 0 0
2
43331 0
0
8 Hex Key~
166 53 87 0 11 12
0 23 22 21 20 0 0 0 0 0
0 48
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
3820 0 0
2
43331 0
0
47
3 1 2 0 0 4224 0 2 11 0 0 5
716 212
792 212
792 237
804 237
804 229
2 2 3 0 0 12416 0 4 2 0 0 5
708 398
708 312
658 312
658 221
671 221
2 1 4 0 0 8320 0 3 2 0 0 5
705 272
705 231
663 231
663 203
671 203
1 0 5 0 0 0 0 3 0 0 6 2
705 308
705 308
1 0 6 0 0 0 0 4 0 0 20 2
708 434
708 434
4 1 5 0 0 4224 0 5 12 0 0 5
646 308
792 308
792 338
804 338
804 330
14 2 7 0 0 12416 0 22 5 0 0 7
507 434
507 477
624 477
624 350
553 350
553 308
601 308
2 3 8 0 0 8320 0 6 5 0 0 4
589 393
593 393
593 317
601 317
2 1 9 0 0 8320 0 7 5 0 0 4
591 234
595 234
595 299
601 299
1 5 10 0 0 4224 0 6 8 0 0 2
553 393
555 393
1 5 11 0 0 4224 0 7 9 0 0 2
555 234
556 234
4 13 12 0 0 4224 0 8 22 0 0 2
505 407
507 407
3 12 13 0 0 4224 0 8 22 0 0 2
505 398
507 398
2 11 14 0 0 4224 0 8 22 0 0 2
505 389
507 389
1 10 15 0 0 4224 0 8 22 0 0 2
505 380
507 380
4 13 16 0 0 4224 0 9 23 0 0 2
506 248
508 248
3 12 17 0 0 4224 0 9 23 0 0 2
506 239
508 239
2 11 18 0 0 4224 0 9 23 0 0 2
506 230
508 230
1 10 19 0 0 4224 0 9 23 0 0 2
506 221
508 221
2 1 6 0 0 4224 0 10 13 0 0 3
621 434
805 434
805 421
14 1 7 0 0 128 0 22 10 0 0 2
507 434
585 434
4 1 20 0 0 8320 0 27 22 0 0 3
44 111
44 353
443 353
3 2 21 0 0 8320 0 27 22 0 0 3
50 111
50 362
443 362
2 3 22 0 0 8320 0 27 22 0 0 3
56 111
56 371
443 371
1 4 23 0 0 8320 0 27 22 0 0 3
62 111
62 380
443 380
14 9 24 0 0 8320 0 23 22 0 0 6
508 275
511 275
511 449
435 449
435 434
443 434
4 1 25 0 0 8320 0 26 23 0 0 3
88 111
88 194
444 194
3 2 26 0 0 8320 0 26 23 0 0 3
94 111
94 203
444 203
2 3 27 0 0 8320 0 26 23 0 0 3
100 111
100 212
444 212
1 4 28 0 0 8320 0 26 23 0 0 5
106 111
106 216
436 216
436 221
444 221
1 9 29 0 0 12416 0 1 23 0 0 6
484 315
517 315
517 290
436 290
436 275
444 275
2 8 30 0 0 8320 0 18 23 0 0 4
360 330
426 330
426 257
444 257
2 7 31 0 0 4224 0 19 23 0 0 4
360 297
431 297
431 248
444 248
2 6 32 0 0 4224 0 20 23 0 0 4
359 264
436 264
436 239
444 239
2 5 33 0 0 4224 0 21 23 0 0 4
359 231
436 231
436 230
444 230
1 1 34 0 0 4224 0 24 18 0 0 3
265 110
265 330
324 330
2 1 35 0 0 4224 0 24 19 0 0 3
259 110
259 297
324 297
3 1 36 0 0 4224 0 24 20 0 0 3
253 110
253 264
323 264
4 1 37 0 0 4224 0 24 21 0 0 3
247 110
247 231
323 231
2 8 38 0 0 8320 0 14 22 0 0 4
360 501
425 501
425 416
443 416
2 7 39 0 0 4224 0 15 22 0 0 4
360 464
430 464
430 407
443 407
2 6 40 0 0 4224 0 16 22 0 0 4
360 428
435 428
435 398
443 398
2 5 41 0 0 4224 0 17 22 0 0 4
360 396
435 396
435 389
443 389
4 1 42 0 0 4224 0 25 17 0 0 3
204 110
204 396
324 396
3 1 43 0 0 4224 0 25 16 0 0 3
210 110
210 428
324 428
2 1 44 0 0 4224 0 25 15 0 0 3
216 110
216 464
324 464
1 1 45 0 0 4224 0 25 14 0 0 3
222 110
222 501
324 501
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
418 541 607 565
428 549 596 565
21 8 BIT COMPARATOR(2'S)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
809 199 854 223
819 207 843 223
3 A>B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
809 298 854 322
819 306 843 322
3 A=B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
220 13 249 37
230 21 238 37
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
62 15 91 39
72 23 80 39
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
811 392 856 416
821 400 845 416
3 A<B
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
