CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
10 10 30 70 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
33
13 Logic Switch~
5 63 353 0 10 11
0 33 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43335 0
0
13 Logic Switch~
5 64 294 0 10 11
0 22 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
43335 0
0
13 Logic Switch~
5 66 239 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
43335 0
0
13 Logic Switch~
5 67 151 0 10 11
0 32 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3421 0 0
2
43335 0
0
13 Logic Switch~
5 69 96 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8157 0 0
2
43335 0
0
13 Logic Switch~
5 70 45 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5572 0 0
2
43335 0
0
14 Logic Display~
6 963 755 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8901 0 0
2
43335 0
0
14 Logic Display~
6 851 755 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7361 0 0
2
43335 0
0
14 Logic Display~
6 643 755 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4747 0 0
2
43335 0
0
14 Logic Display~
6 433 755 0 1 2
10 25
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
972 0 0
2
43335 0
0
14 Logic Display~
6 260 754 0 1 2
10 34
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3472 0 0
2
43335 0
0
14 Logic Display~
6 145 755 0 1 2
10 37
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9998 0 0
2
43335 0
0
8 2-In OR~
219 873 506 0 3 22
0 4 3 2
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
3536 0 0
2
43335 0
0
9 2-In AND~
219 789 394 0 3 22
0 10 11 8
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U11A
-15 -11 13 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
4597 0 0
2
43335 0
0
8 2-In OR~
219 665 511 0 3 22
0 13 12 9
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3835 0 0
2
43335 0
0
9 2-In AND~
219 587 394 0 3 22
0 11 21 15
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3D
-12 -11 9 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
3670 0 0
2
43335 0
0
9 2-In AND~
219 549 395 0 3 22
0 22 10 17
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3C
-12 -11 9 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
5616 0 0
2
43335 0
0
8 2-In OR~
219 441 513 0 3 22
0 24 23 20
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
9323 0 0
2
43335 0
0
9 2-In AND~
219 398 396 0 3 22
0 11 32 26
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3B
-12 -11 9 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
317 0 0
2
43335 0
0
9 2-In AND~
219 358 396 0 3 22
0 22 21 31
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3A
-12 -11 9 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3108 0 0
2
43335 0
0
9 2-In AND~
219 317 397 0 3 22
0 33 10 30
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1D
-12 -11 9 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
4299 0 0
2
43335 0
0
9 2-In AND~
219 213 396 0 3 22
0 22 32 35
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1C
-12 -11 9 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
9672 0 0
2
43335 0
0
9 2-In AND~
219 169 396 0 3 22
0 33 21 36
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1B
-12 -10 9 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
7876 0 0
2
43335 0
0
9 2-In AND~
219 121 397 0 3 22
0 32 33 37
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1A
-12 -10 9 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
6369 0 0
2
43335 0
0
2 HA
94 190 471 0 4 9
0 35 36 28 34
2 HA
1 0 656 0
0
2 U2
-7 -28 7 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 U
9172 0 0
2
43334.7 0
0
2 HA
94 355 469 0 4 9
0 31 30 24 29
2 HA
2 0 656 0
0
2 U4
-7 -28 7 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 U
7100 0 0
2
43334.7 0
0
2 HA
94 354 554 0 4 9
0 28 29 23 27
2 HA
3 0 656 0
0
2 U5
-7 -28 7 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 U
3820 0 0
2
43334.7 0
0
2 HA
94 354 637 0 4 9
0 26 27 19 25
2 HA
4 0 656 0
0
2 U6
-7 -28 7 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 U
7678 0 0
2
43334.7 0
0
2 HA
94 568 465 0 4 9
0 19 20 13 18
2 HA
5 0 656 0
0
2 U8
-7 -28 7 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 U
961 0 0
2
43334.7 0
0
2 HA
94 569 552 0 4 9
0 17 18 12 16
2 HA
6 0 656 0
0
2 U9
-7 -28 7 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 U
3178 0 0
2
43334.7 0
0
2 HA
94 568 635 0 4 9
0 15 16 7 14
2 HA
7 0 656 0
0
3 U10
-11 -28 10 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 U
3409 0 0
2
43334.7 0
0
2 HA
94 787 460 0 4 9
0 8 9 4 6
2 HA
8 0 656 0
0
3 U12
-11 -28 10 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 U
3951 0 0
2
43334.7 0
0
2 HA
94 786 548 0 4 9
0 6 7 3 5
2 HA
9 0 656 0
0
3 U13
-11 -28 10 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 U
8885 0 0
2
43334.7 0
0
54
3 1 2 0 0 8320 0 13 7 0 0 7
906 506
947 506
947 774
951 774
951 781
963 781
963 773
3 2 3 0 0 8320 0 33 13 0 0 4
819 557
852 557
852 515
860 515
3 1 4 0 0 4224 0 32 13 0 0 4
820 469
852 469
852 497
860 497
4 1 5 0 0 8320 0 33 8 0 0 7
819 548
834 548
834 773
839 773
839 781
851 781
851 773
4 1 6 0 0 12416 0 32 33 0 0 6
820 460
833 460
833 503
729 503
729 548
753 548
3 2 7 0 0 4224 0 31 33 0 0 4
601 644
745 644
745 557
753 557
3 1 8 0 0 4224 0 14 32 0 0 4
787 417
737 417
737 460
754 460
3 2 9 0 0 4224 0 15 32 0 0 4
698 511
746 511
746 469
754 469
1 0 10 0 0 4096 0 14 0 0 54 2
796 372
796 45
2 0 11 0 0 4096 0 14 0 0 51 2
778 372
778 239
3 2 12 0 0 4224 0 30 15 0 0 4
602 561
644 561
644 520
652 520
3 1 13 0 0 4224 0 29 15 0 0 4
601 474
644 474
644 502
652 502
4 1 14 0 0 8320 0 31 9 0 0 7
601 635
625 635
625 773
631 773
631 781
643 781
643 773
3 1 15 0 0 8320 0 16 31 0 0 6
585 417
617 417
617 601
513 601
513 635
535 635
4 2 16 0 0 12416 0 30 31 0 0 6
602 552
625 552
625 592
503 592
503 644
535 644
3 1 17 0 0 8320 0 17 30 0 0 4
547 418
518 418
518 552
536 552
4 2 18 0 0 12416 0 29 30 0 0 6
601 465
625 465
625 503
510 503
510 561
536 561
3 1 19 0 0 8320 0 28 29 0 0 4
387 646
486 646
486 465
535 465
3 2 20 0 0 4224 0 18 29 0 0 4
474 513
527 513
527 474
535 474
1 0 11 0 0 0 0 16 0 0 51 2
594 372
594 239
2 0 21 0 0 4096 0 16 0 0 53 2
576 372
576 96
1 0 22 0 0 4096 0 17 0 0 50 2
556 373
556 294
2 0 10 0 0 4096 0 17 0 0 54 2
538 373
538 45
3 2 23 0 0 8320 0 27 18 0 0 4
387 563
420 563
420 522
428 522
3 1 24 0 0 4224 0 26 18 0 0 4
388 478
420 478
420 504
428 504
4 1 25 0 0 8320 0 28 10 0 0 7
387 637
412 637
412 773
421 773
421 781
433 781
433 773
3 1 26 0 0 4224 0 19 28 0 0 5
396 419
396 601
276 601
276 637
321 637
4 2 27 0 0 12416 0 27 28 0 0 6
387 554
412 554
412 592
285 592
285 646
321 646
3 1 28 0 0 8320 0 25 27 0 0 4
223 480
284 480
284 554
321 554
4 2 29 0 0 12416 0 26 27 0 0 6
388 469
411 469
411 512
292 512
292 563
321 563
3 2 30 0 0 12416 0 21 26 0 0 5
315 420
315 427
293 427
293 478
322 478
3 1 31 0 0 8320 0 20 26 0 0 5
356 419
356 433
299 433
299 469
322 469
1 0 11 0 0 4096 0 19 0 0 51 2
405 374
405 239
2 0 32 0 0 4096 0 19 0 0 52 2
387 374
387 151
1 0 22 0 0 4096 0 20 0 0 50 2
365 374
365 294
2 0 21 0 0 4096 0 20 0 0 53 2
347 374
347 96
1 0 33 0 0 4096 0 21 0 0 49 2
324 375
324 353
2 0 10 0 0 4096 0 21 0 0 54 2
306 375
306 45
4 1 34 0 0 8320 0 25 11 0 0 7
223 471
236 471
236 773
248 773
248 780
260 780
260 772
3 1 35 0 0 8320 0 22 25 0 0 5
211 419
211 428
143 428
143 471
157 471
3 2 36 0 0 8320 0 23 25 0 0 4
167 419
134 419
134 480
157 480
1 0 22 0 0 0 0 22 0 0 50 2
220 374
220 294
2 0 32 0 0 0 0 22 0 0 52 2
202 374
202 151
1 0 33 0 0 0 0 23 0 0 49 2
176 374
176 353
2 0 21 0 0 0 0 23 0 0 53 2
158 374
158 96
3 1 37 0 0 4224 0 24 12 0 0 6
119 420
119 773
133 773
133 781
145 781
145 773
1 0 32 0 0 4096 0 24 0 0 52 2
128 375
128 151
2 0 33 0 0 0 0 24 0 0 49 2
110 375
110 353
1 0 33 0 0 4224 0 1 0 0 0 2
75 353
1156 353
1 0 22 0 0 4224 0 2 0 0 0 2
76 294
1155 294
1 0 11 0 0 4224 0 3 0 0 0 2
78 239
1156 239
1 0 32 0 0 4224 0 4 0 0 0 2
79 151
1156 151
1 0 21 0 0 4224 0 5 0 0 0 2
81 96
1155 96
1 0 10 0 0 4224 0 6 0 0 0 2
82 45
1155 45
12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
944 702 981 726
954 710 970 726
2 S5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
833 704 870 728
843 712 859 728
2 S4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
624 705 661 729
634 713 650 729
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
415 703 452 727
425 711 441 727
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
242 702 279 726
252 710 268 726
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
127 702 164 726
137 710 153 726
2 SO
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
16 329 53 353
26 337 42 353
2 B0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
17 273 54 297
27 281 43 297
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
18 215 55 239
28 223 44 239
2 B2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
19 127 56 151
29 135 45 151
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
20 74 57 98
30 82 46 98
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
20 23 57 47
30 31 46 47
2 A2
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
