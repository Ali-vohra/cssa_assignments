CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
14
13 Logic Switch~
5 414 310 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V4
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4900 0 0
2
5.89862e-315 0
0
13 Logic Switch~
5 302 309 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V3
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8783 0 0
2
5.89862e-315 0
0
13 Logic Switch~
5 197 310 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V2
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3221 0 0
2
5.89862e-315 0
0
13 Logic Switch~
5 125 123 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3215 0 0
2
5.89862e-315 0
0
5 4082~
219 485 194 0 5 22
0 7 4 3 2 8
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U3B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 3 0
1 U
7903 0 0
2
5.89862e-315 0
0
5 4082~
219 486 144 0 5 22
0 7 4 5 2 9
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U3A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 3 0
1 U
7121 0 0
2
5.89862e-315 0
0
5 4082~
219 487 96 0 5 22
0 7 6 3 2 10
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U2B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 2 0
1 U
4484 0 0
2
5.89862e-315 0
0
5 4082~
219 488 47 0 5 22
0 7 6 5 2 11
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U2A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 2 0
1 U
5996 0 0
2
5.89862e-315 0
0
9 Inverter~
13 393 259 0 2 22
0 6 4
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U1B
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
7804 0 0
2
5.89862e-315 0
0
9 Inverter~
13 281 260 0 2 22
0 5 3
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U1A
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
5523 0 0
2
5.89862e-315 0
0
14 Logic Display~
6 641 183 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3330 0 0
2
5.89862e-315 0
0
14 Logic Display~
6 642 128 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3465 0 0
2
5.89862e-315 0
0
14 Logic Display~
6 641 78 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8396 0 0
2
5.89862e-315 0
0
14 Logic Display~
6 641 25 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3685 0 0
2
5.89862e-315 0
0
27
4 0 2 0 0 4096 0 5 0 0 23 2
461 208
198 208
4 0 2 0 0 4096 0 6 0 0 23 2
462 158
198 158
4 0 2 0 0 4096 0 7 0 0 23 2
463 110
198 110
3 0 3 0 0 4096 0 5 0 0 18 2
461 199
284 199
2 0 4 0 0 4096 0 5 0 0 17 2
461 190
396 190
3 0 5 0 0 4096 0 6 0 0 22 2
462 149
303 149
2 0 4 0 0 4096 0 6 0 0 17 2
462 140
396 140
3 0 3 0 0 4096 0 7 0 0 18 2
463 101
284 101
2 0 6 0 0 4096 0 7 0 0 21 2
463 92
415 92
4 0 2 0 0 4096 0 8 0 0 23 2
464 61
198 61
3 0 5 0 0 4096 0 8 0 0 22 2
464 52
303 52
2 0 6 0 0 4096 0 8 0 0 21 2
464 43
415 43
1 1 7 0 0 4096 0 5 4 0 0 4
461 181
161 181
161 123
137 123
1 1 7 0 0 4096 0 6 4 0 0 4
462 131
156 131
156 123
137 123
1 1 7 0 0 4096 0 7 4 0 0 4
463 83
151 83
151 123
137 123
1 1 7 0 0 4224 0 8 4 0 0 4
464 34
146 34
146 123
137 123
2 0 4 0 0 4224 0 9 0 0 0 2
396 241
396 14
2 0 3 0 0 4224 0 10 0 0 0 2
284 242
284 14
1 1 5 0 0 0 0 2 10 0 0 4
303 296
303 286
284 286
284 278
1 1 6 0 0 0 0 1 9 0 0 4
415 297
415 285
396 285
396 277
1 0 6 0 0 4224 0 1 0 0 0 2
415 297
415 14
1 0 5 0 0 4224 0 2 0 0 0 2
303 296
303 13
1 0 2 0 0 4224 0 3 0 0 0 2
198 297
198 12
5 1 8 0 0 4224 0 5 11 0 0 5
506 194
629 194
629 209
641 209
641 201
5 1 9 0 0 4224 0 6 12 0 0 5
507 144
630 144
630 154
642 154
642 146
5 1 10 0 0 4224 0 7 13 0 0 5
508 96
629 96
629 104
641 104
641 96
5 1 11 0 0 4224 0 8 14 0 0 3
509 47
641 47
641 43
8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
70 100 107 124
80 108 96 124
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
661 9 698 33
671 17 687 33
2 D3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
663 62 700 86
673 70 689 86
2 D2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
665 113 702 137
675 121 691 137
2 D1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
665 169 702 193
675 177 691 193
2 D0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
184 328 213 352
194 336 202 352
1 E
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
398 329 435 353
408 337 424 353
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
284 329 321 353
294 337 310 353
2 S0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
