CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
16
13 Logic Switch~
5 745 560 0 1 11
0 6
0
0 0 21360 90
2 0V
14 0 28 8
3 V11
10 -10 31 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43361.9 0
0
13 Logic Switch~
5 646 561 0 1 11
0 7
0
0 0 21360 90
2 0V
14 0 28 8
3 V10
10 -10 31 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
43361.9 0
0
13 Logic Switch~
5 560 560 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V9
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
43361.9 0
0
13 Logic Switch~
5 103 480 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3421 0 0
2
43361.9 0
0
13 Logic Switch~
5 104 416 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8157 0 0
2
43361.9 0
0
13 Logic Switch~
5 105 354 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5572 0 0
2
43361.9 0
0
13 Logic Switch~
5 105 293 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8901 0 0
2
43361.9 0
0
13 Logic Switch~
5 105 234 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7361 0 0
2
43361.9 0
0
13 Logic Switch~
5 106 179 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4747 0 0
2
43361.9 0
0
13 Logic Switch~
5 107 125 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
972 0 0
2
43361.9 0
0
13 Logic Switch~
5 107 74 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3472 0 0
2
43361.9 0
0
14 Logic Display~
6 977 264 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9998 0 0
2
43361.9 0
0
8 2-In OR~
219 840 278 0 3 22
0 4 3 2
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3536 0 0
2
43361.9 0
0
9 Inverter~
13 533 508 0 2 22
0 8 5
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U3A
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
4597 0 0
2
43361.9 0
0
8 4x1 MUX~
94 430 155 0 8 17
0 16 15 14 13 4 7 6 5
7 4x1 MUX
1 0 560 0
0
2 U1
1 -68 15 -60
0
0
0
0
0
0
17

0 3 4 5 6 9 12 13 16 3
4 5 6 9 12 13 16 0
0 0 0 0 0 0 0 0
1 U
3835 0 0
2
43361.9 0
0
8 4x1 MUX~
94 427 374 0 8 17
0 12 11 10 9 3 7 6 8
7 4x1 MUX
2 0 560 0
0
2 U2
1 -68 15 -60
0
0
0
0
0
0
17

0 3 4 5 6 9 12 13 16 3
4 5 6 9 12 13 16 0
0 0 0 0 0 0 0 0
1 U
3670 0 0
2
43361.9 0
0
18
3 1 2 0 0 4224 0 13 12 0 0 5
873 278
965 278
965 290
977 290
977 282
5 2 3 0 0 4224 0 16 13 0 0 4
476 420
819 420
819 287
827 287
5 1 4 0 0 4224 0 15 13 0 0 4
479 201
819 201
819 269
827 269
8 2 5 0 0 8320 0 15 14 0 0 3
479 120
536 120
536 490
1 7 6 0 0 8192 0 1 16 0 0 3
746 547
746 374
476 374
1 7 6 0 0 4224 0 1 15 0 0 3
746 547
746 155
479 155
1 6 7 0 0 8192 0 2 16 0 0 3
647 548
647 385
476 385
1 6 7 0 0 4224 0 2 15 0 0 3
647 548
647 166
479 166
1 8 8 0 0 4224 0 3 16 0 0 3
561 547
561 339
476 339
1 1 8 0 0 0 0 3 14 0 0 4
561 547
561 534
536 534
536 526
1 4 9 0 0 4224 0 4 16 0 0 4
115 480
381 480
381 397
394 397
1 3 10 0 0 4224 0 5 16 0 0 4
116 416
386 416
386 385
394 385
1 2 11 0 0 4224 0 6 16 0 0 4
117 354
381 354
381 374
394 374
1 1 12 0 0 4224 0 7 16 0 0 4
117 293
386 293
386 363
394 363
1 4 13 0 0 4224 0 8 15 0 0 4
117 234
384 234
384 178
397 178
1 3 14 0 0 4224 0 9 15 0 0 4
118 179
389 179
389 166
397 166
1 2 15 0 0 4224 0 10 15 0 0 4
119 125
384 125
384 155
397 155
1 1 16 0 0 4224 0 11 15 0 0 4
119 74
389 74
389 144
397 144
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
