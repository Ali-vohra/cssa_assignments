CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 60 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
45
13 Logic Switch~
5 63 545 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 60 401 0 10 11
0 50 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
43335 0
0
13 Logic Switch~
5 60 351 0 10 11
0 48 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3124 0 0
2
43335 1
0
13 Logic Switch~
5 60 302 0 10 11
0 46 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
43335 2
0
13 Logic Switch~
5 60 254 0 10 11
0 44 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8157 0 0
2
43335 3
0
13 Logic Switch~
5 57 167 0 10 11
0 49 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5572 0 0
2
43335 4
0
13 Logic Switch~
5 57 121 0 10 11
0 47 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8901 0 0
2
43335 5
0
13 Logic Switch~
5 57 73 0 10 11
0 45 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7361 0 0
2
43335 6
0
13 Logic Switch~
5 58 32 0 10 11
0 43 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4747 0 0
2
43335 7
0
14 Logic Display~
6 1532 923 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
972 0 0
2
43335 0
0
14 Logic Display~
6 1417 930 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3472 0 0
2
43335 0
0
14 Logic Display~
6 1260 930 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9998 0 0
2
43335 0
0
14 Logic Display~
6 1045 935 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3536 0 0
2
43335 0
0
14 Logic Display~
6 798 933 0 1 2
10 24
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4597 0 0
2
43335 0
0
14 Logic Display~
6 532 933 0 1 2
10 33
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3835 0 0
2
43335 0
0
14 Logic Display~
6 312 935 0 1 2
10 39
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3670 0 0
2
43335 0
0
14 Logic Display~
6 170 938 0 1 2
10 42
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5616 0 0
2
43335 0
0
9 2-In AND~
219 1302 444 0 3 22
0 43 44 4
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U14D
-14 -10 14 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
9323 0 0
2
43335 8
0
9 2-In AND~
219 1125 445 0 3 22
0 44 45 8
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U14C
-15 -11 13 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
317 0 0
2
43335 9
0
9 2-In AND~
219 1083 446 0 3 22
0 46 43 9
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U14B
-15 -10 13 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3108 0 0
2
43335 10
0
9 2-In AND~
219 907 445 0 3 22
0 44 47 18
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U14A
-15 -10 13 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
4299 0 0
2
43335 11
0
9 2-In AND~
219 866 446 0 3 22
0 46 45 19
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U8D
-12 -10 9 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
9672 0 0
2
43335 12
0
9 2-In AND~
219 826 446 0 3 22
0 48 43 20
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U8C
-12 -9 9 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
7876 0 0
2
43335 13
0
9 2-In AND~
219 654 447 0 3 22
0 44 49 27
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U8B
-12 -9 9 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
6369 0 0
2
43335 14
0
9 2-In AND~
219 614 447 0 3 22
0 46 47 28
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U8A
-12 -9 9 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
9172 0 0
2
43335 15
0
9 2-In AND~
219 572 448 0 3 22
0 48 45 29
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3D
-11 -9 10 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
7100 0 0
2
43335 16
0
9 2-In AND~
219 530 449 0 3 22
0 50 43 30
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3C
-11 -8 10 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
3820 0 0
2
43335 17
0
9 2-In AND~
219 366 450 0 3 22
0 46 49 36
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3B
-12 -9 9 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
7678 0 0
2
43335 18
0
9 2-In AND~
219 320 451 0 3 22
0 48 47 37
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3A
-12 -9 9 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
961 0 0
2
43335 19
0
9 2-In AND~
219 275 451 0 3 22
0 50 45 38
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1D
-12 -8 9 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
3178 0 0
2
43335 20
0
9 2-In AND~
219 207 450 0 3 22
0 48 49 40
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1C
-12 -6 9 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3409 0 0
2
43335 21
0
9 2-In AND~
219 158 451 0 3 22
0 50 47 41
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1B
-12 -6 9 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3951 0 0
2
43335 22
0
9 2-In AND~
219 108 450 0 3 22
0 50 49 42
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1A
-12 -5 9 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
8885 0 0
2
43335 23
0
2 FA
94 182 531 0 5 11
0 41 40 15 34 39
2 FA
1 0 688 0
0
2 U2
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 1 0 0 0
1 U
3780 0 0
2
5.89859e-315 0
0
2 FA
94 321 530 0 5 11
0 36 37 38 32 35
2 FA
2 0 688 0
0
2 U4
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 1 0 0 0
1 U
9265 0 0
2
5.89859e-315 0
0
2 FA
94 319 619 0 5 11
0 34 35 15 31 33
2 FA
3 0 688 0
0
2 U5
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
9442 0 0
2
43334.9 0
0
2 FA
94 595 530 0 5 11
0 30 31 32 23 26
2 FA
4 0 688 0
0
2 U6
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
9424 0 0
2
43334.9 0
0
2 FA
94 595 616 0 5 11
0 27 28 29 22 25
2 FA
5 0 688 0
0
2 U7
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
9968 0 0
2
43334.9 0
0
2 FA
94 596 713 0 5 11
0 25 26 15 21 24
2 FA
6 0 688 0
0
2 U9
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
9281 0 0
2
43334.9 0
0
2 FA
94 866 525 0 5 11
0 23 22 21 13 17
2 FA
7 0 688 0
0
3 U10
-11 -29 10 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
8464 0 0
2
43334.9 0
0
2 FA
94 867 611 0 5 11
0 18 19 20 12 16
2 FA
8 0 688 0
0
3 U11
-11 -29 10 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
7168 0 0
2
43334.9 0
0
2 FA
94 865 708 0 5 11
0 16 17 15 11 14
2 FA
9 0 688 0
0
3 U12
-11 -29 10 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
3171 0 0
2
43334.9 0
0
2 FA
94 1105 522 0 5 11
0 13 12 11 6 10
2 FA
10 0 688 0
0
3 U13
-11 -29 10 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
4139 0 0
2
43334.9 0
0
2 FA
94 1105 606 0 5 11
0 8 9 10 5 7
2 FA
11 0 688 0
0
3 U15
-11 -29 10 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
6435 0 0
2
43334.9 0
0
2 FA
94 1301 519 0 5 11
0 6 5 4 2 3
2 FA
12 0 688 0
0
3 U16
-11 -29 10 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
5283 0 0
2
43334.9 0
0
84
4 1 2 0 0 8320 0 45 10 0 0 5
1334 537
1468 537
1468 961
1532 961
1532 941
5 1 3 0 0 8320 0 45 11 0 0 5
1334 519
1357 519
1357 962
1417 962
1417 948
3 3 4 0 0 8320 0 18 45 0 0 4
1300 467
1255 467
1255 537
1268 537
4 2 5 0 0 8320 0 44 45 0 0 4
1138 624
1200 624
1200 528
1268 528
4 1 6 0 0 12416 0 43 45 0 0 4
1138 540
1189 540
1189 519
1268 519
5 1 7 0 0 8320 0 44 12 0 0 5
1138 606
1155 606
1155 962
1260 962
1260 948
3 1 8 0 0 12416 0 19 44 0 0 5
1123 468
1123 486
1034 486
1034 606
1072 606
3 2 9 0 0 12416 0 20 44 0 0 5
1081 469
1081 477
1044 477
1044 615
1072 615
5 3 10 0 0 12416 0 43 44 0 0 6
1138 522
1155 522
1155 567
1053 567
1053 624
1072 624
4 3 11 0 0 8320 0 42 43 0 0 4
898 726
950 726
950 540
1072 540
4 2 12 0 0 12416 0 41 43 0 0 4
900 629
939 629
939 531
1072 531
4 1 13 0 0 12416 0 40 43 0 0 4
899 543
929 543
929 522
1072 522
5 1 14 0 0 8320 0 42 13 0 0 5
898 708
921 708
921 963
1045 963
1045 953
0 3 15 0 0 8320 0 0 42 34 0 5
152 637
152 677
799 677
799 726
832 726
5 1 16 0 0 12416 0 41 42 0 0 6
900 611
914 611
914 663
814 663
814 708
832 708
5 2 17 0 0 8320 0 40 42 0 0 6
899 525
921 525
921 656
808 656
808 717
832 717
3 1 18 0 0 12416 0 21 41 0 0 5
905 468
905 485
808 485
808 611
834 611
3 2 19 0 0 12416 0 22 41 0 0 5
864 469
864 477
816 477
816 620
834 620
3 3 20 0 0 4224 0 23 41 0 0 3
824 469
824 629
834 629
4 3 21 0 0 8320 0 39 40 0 0 4
629 731
682 731
682 543
833 543
4 2 22 0 0 12416 0 38 40 0 0 4
628 634
674 634
674 534
833 534
4 1 23 0 0 8320 0 37 40 0 0 3
628 548
628 525
833 525
5 1 24 0 0 8320 0 39 14 0 0 5
629 713
667 713
667 963
798 963
798 951
0 3 15 0 0 0 0 0 39 34 0 3
84 637
84 731
563 731
5 1 25 0 0 12416 0 38 39 0 0 6
628 616
662 616
662 667
519 667
519 713
563 713
5 2 26 0 0 12416 0 37 39 0 0 6
628 530
668 530
668 662
513 662
513 722
563 722
3 1 27 0 0 8320 0 24 38 0 0 5
652 470
652 497
504 497
504 616
562 616
3 2 28 0 0 12416 0 25 38 0 0 5
612 470
612 490
512 490
512 625
562 625
3 3 29 0 0 12416 0 26 38 0 0 5
570 471
570 483
520 483
520 634
562 634
3 1 30 0 0 4224 0 27 37 0 0 3
528 472
528 530
562 530
4 2 31 0 0 12416 0 36 37 0 0 4
352 637
399 637
399 539
562 539
4 3 32 0 0 4224 0 35 37 0 0 2
354 548
562 548
5 1 33 0 0 8320 0 36 15 0 0 5
352 619
379 619
379 964
532 964
532 951
1 3 15 0 0 0 0 1 36 0 0 3
75 545
75 637
286 637
4 1 34 0 0 8320 0 34 36 0 0 3
215 549
215 619
286 619
5 2 35 0 0 12416 0 35 36 0 0 6
354 530
379 530
379 576
257 576
257 628
286 628
3 1 36 0 0 8320 0 28 35 0 0 5
364 473
364 486
258 486
258 530
288 530
3 2 37 0 0 8320 0 29 35 0 0 5
318 474
318 493
266 493
266 539
288 539
3 3 38 0 0 4224 0 30 35 0 0 3
273 474
273 548
288 548
1 3 15 0 0 128 0 1 34 0 0 3
75 545
75 549
149 549
5 1 39 0 0 8320 0 34 16 0 0 5
215 531
235 531
235 963
312 963
312 953
3 2 40 0 0 8320 0 31 34 0 0 5
205 473
205 488
136 488
136 540
149 540
3 1 41 0 0 8320 0 32 34 0 0 4
156 474
121 474
121 531
149 531
3 1 42 0 0 4224 0 33 17 0 0 4
106 473
106 962
170 962
170 956
1 0 43 0 0 4096 0 18 0 0 84 2
1309 422
1309 32
2 0 44 0 0 4096 0 18 0 0 80 2
1291 422
1291 254
1 0 44 0 0 4096 0 19 0 0 80 2
1132 423
1132 254
2 0 45 0 0 4096 0 19 0 0 83 2
1114 423
1114 73
1 0 46 0 0 4096 0 20 0 0 79 2
1090 424
1090 302
2 0 43 0 0 4096 0 20 0 0 84 2
1072 424
1072 32
1 0 44 0 0 0 0 21 0 0 80 2
914 423
914 254
2 0 47 0 0 4096 0 21 0 0 82 2
896 423
896 121
1 0 46 0 0 0 0 22 0 0 79 2
873 424
873 302
2 0 45 0 0 4096 0 22 0 0 83 2
855 424
855 73
1 0 48 0 0 4096 0 23 0 0 78 2
833 424
833 351
2 0 43 0 0 0 0 23 0 0 84 2
815 424
815 32
1 0 44 0 0 4096 0 24 0 0 80 2
661 425
661 254
2 0 49 0 0 4096 0 24 0 0 81 2
643 425
643 167
1 0 46 0 0 4096 0 25 0 0 79 2
621 425
621 302
2 0 47 0 0 4096 0 25 0 0 82 2
603 425
603 121
1 0 48 0 0 4096 0 26 0 0 78 2
579 426
579 351
2 0 45 0 0 4096 0 26 0 0 83 2
561 426
561 73
1 0 50 0 0 4096 0 27 0 0 77 2
537 427
537 401
2 0 43 0 0 4096 0 27 0 0 84 2
519 427
519 32
1 0 46 0 0 4096 0 28 0 0 79 2
373 428
373 302
2 0 49 0 0 4096 0 28 0 0 81 2
355 428
355 167
1 0 48 0 0 4096 0 29 0 0 78 2
327 429
327 351
2 0 47 0 0 4096 0 29 0 0 82 2
309 429
309 121
1 0 50 0 0 4096 0 30 0 0 77 2
282 429
282 401
2 0 45 0 0 4096 0 30 0 0 83 2
264 429
264 73
1 0 48 0 0 0 0 31 0 0 78 2
214 428
214 351
2 0 49 0 0 0 0 31 0 0 81 2
196 428
196 167
1 0 50 0 0 0 0 32 0 0 77 2
165 429
165 401
2 0 47 0 0 0 0 32 0 0 82 2
147 429
147 121
2 0 49 0 0 0 0 33 0 0 81 2
97 428
97 167
1 0 50 0 0 0 0 33 0 0 77 2
115 428
115 401
1 0 50 0 0 4224 0 2 0 0 0 2
72 401
1552 401
1 0 48 0 0 4224 0 3 0 0 0 2
72 351
1552 351
1 0 46 0 0 4224 0 4 0 0 0 2
72 302
1551 302
1 0 44 0 0 4224 0 5 0 0 0 2
72 254
1551 254
1 0 49 0 0 4224 0 6 0 0 0 2
69 167
1551 167
1 0 47 0 0 4224 0 7 0 0 0 2
69 121
1551 121
1 0 45 0 0 4224 0 8 0 0 0 2
69 73
1552 73
1 0 43 0 0 4224 0 9 0 0 0 2
70 32
1552 32
16
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1507 866 1559 885
1524 879 1541 892
2 S7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1391 868 1443 887
1408 881 1425 894
2 S6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1234 867 1286 886
1251 880 1268 893
2 S5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1020 870 1072 889
1037 883 1054 896
2 S4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
773 871 825 890
790 885 807 898
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
507 872 557 891
523 885 540 898
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
286 872 338 891
303 885 320 898
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
146 872 196 891
162 885 179 898
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
10 377 47 401
20 385 36 401
2 B0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
10 332 47 356
20 340 36 356
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
12 283 49 307
22 291 38 307
2 B2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
11 230 48 254
21 238 37 254
2 B3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
8 144 45 168
18 152 34 168
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
8 99 45 123
18 107 34 123
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
7 51 44 75
17 59 33 75
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
7 10 44 34
17 18 33 34
2 A3
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
