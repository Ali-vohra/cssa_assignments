CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
20
13 Logic Switch~
5 567 242 0 1 11
0 6
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 329 277 0 1 11
0 17
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 147 442 0 1 11
0 30
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 152 229 0 10 11
0 31 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
5.89855e-315 0
0
12 Hex Display~
7 782 158 0 18 19
10 2 3 4 5 0 0 0 0 0
0 1 1 1 1 1 1 1 8
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
8157 0 0
2
5.89855e-315 0
0
9 Inverter~
13 472 406 0 2 22
0 7 8
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
5572 0 0
2
5.89855e-315 0
0
5 4030~
219 565 529 0 3 22
0 13 8 9
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U6D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 2 0
1 U
8901 0 0
2
5.89855e-315 0
0
5 4030~
219 564 475 0 3 22
0 14 8 10
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U6C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
7361 0 0
2
5.89855e-315 0
0
5 4030~
219 564 425 0 3 22
0 15 8 11
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U6B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
4747 0 0
2
5.89855e-315 0
0
5 4030~
219 564 374 0 3 22
0 16 8 12
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U6A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
972 0 0
2
5.89855e-315 0
0
6 74LS83
105 669 281 0 14 29
0 6 6 6 6 12 11 10 9 7
5 4 3 2 40
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U5
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
3472 0 0
2
5.89855e-315 0
0
9 Inverter~
13 348 439 0 2 22
0 26 22
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
9998 0 0
2
5.89855e-315 0
0
9 Inverter~
13 347 402 0 2 22
0 27 23
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3536 0 0
2
5.89855e-315 0
0
9 Inverter~
13 347 363 0 2 22
0 28 24
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
4597 0 0
2
5.89855e-315 0
0
9 Inverter~
13 347 326 0 2 22
0 29 25
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3835 0 0
2
5.89855e-315 0
0
6 74LS83
105 460 286 0 14 29
0 21 20 19 18 25 24 23 22 17
16 15 14 13 7
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U3
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
3670 0 0
2
5.89855e-315 0
0
8 Hex Key~
166 156 311 0 11 12
0 32 33 34 35 0 0 0 0 0
9 57
0
0 0 4640 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
5616 0 0
2
5.89855e-315 0
0
8 Hex Key~
166 154 81 0 11 12
0 36 37 38 39 0 0 0 0 0
1 49
0
0 0 4640 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
9323 0 0
2
5.89855e-315 0
0
6 74LS83
105 240 404 0 14 29
0 35 34 33 32 30 30 31 30 30
29 28 27 26 41
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U2
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
317 0 0
2
5.89855e-315 0
0
6 74LS83
105 241 200 0 14 29
0 39 38 37 36 30 30 31 30 30
21 20 19 18 42
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
3108 0 0
2
5.89855e-315 0
0
53
13 1 2 0 0 8320 0 11 5 0 0 3
701 299
791 299
791 182
12 2 3 0 0 8320 0 11 5 0 0 3
701 290
785 290
785 182
11 3 4 0 0 8320 0 11 5 0 0 3
701 281
779 281
779 182
10 4 5 0 0 8320 0 11 5 0 0 3
701 272
773 272
773 182
1 4 6 0 0 4096 0 1 11 0 0 4
579 242
614 242
614 272
637 272
1 3 6 0 0 4096 0 1 11 0 0 4
579 242
619 242
619 263
637 263
1 2 6 0 0 4096 0 1 11 0 0 4
579 242
624 242
624 254
637 254
1 1 6 0 0 4224 0 1 11 0 0 4
579 242
629 242
629 245
637 245
14 9 7 0 0 4224 0 16 11 0 0 4
492 331
609 331
609 326
637 326
2 2 8 0 0 8320 0 6 7 0 0 4
493 406
511 406
511 538
549 538
2 2 8 0 0 0 0 6 8 0 0 4
493 406
515 406
515 484
548 484
2 2 8 0 0 0 0 6 9 0 0 4
493 406
520 406
520 434
548 434
2 2 8 0 0 0 0 6 10 0 0 4
493 406
540 406
540 383
548 383
14 1 7 0 0 0 0 16 6 0 0 6
492 331
497 331
497 421
449 421
449 406
457 406
3 8 9 0 0 8320 0 7 11 0 0 4
598 529
614 529
614 308
637 308
3 7 10 0 0 8320 0 8 11 0 0 4
597 475
619 475
619 299
637 299
3 6 11 0 0 8320 0 9 11 0 0 4
597 425
624 425
624 290
637 290
3 5 12 0 0 8320 0 10 11 0 0 4
597 374
629 374
629 281
637 281
13 1 13 0 0 8320 0 16 7 0 0 4
492 304
526 304
526 520
549 520
12 1 14 0 0 8320 0 16 8 0 0 4
492 295
530 295
530 466
548 466
11 1 15 0 0 8320 0 16 9 0 0 4
492 286
535 286
535 416
548 416
10 1 16 0 0 8320 0 16 10 0 0 4
492 277
540 277
540 365
548 365
1 9 17 0 0 4224 0 2 16 0 0 4
341 277
400 277
400 331
428 331
13 4 18 0 0 4224 0 20 16 0 0 4
273 218
405 218
405 277
428 277
12 3 19 0 0 4224 0 20 16 0 0 4
273 209
410 209
410 268
428 268
11 2 20 0 0 4224 0 20 16 0 0 4
273 200
415 200
415 259
428 259
10 1 21 0 0 4224 0 20 16 0 0 4
273 191
420 191
420 250
428 250
2 8 22 0 0 8320 0 12 16 0 0 4
369 439
405 439
405 313
428 313
2 7 23 0 0 8320 0 13 16 0 0 4
368 402
410 402
410 304
428 304
2 6 24 0 0 8320 0 14 16 0 0 4
368 363
415 363
415 295
428 295
2 5 25 0 0 4224 0 15 16 0 0 4
368 326
420 326
420 286
428 286
13 1 26 0 0 4224 0 19 12 0 0 4
272 422
325 422
325 439
333 439
12 1 27 0 0 4224 0 19 13 0 0 4
272 413
324 413
324 402
332 402
11 1 28 0 0 4224 0 19 14 0 0 4
272 404
319 404
319 363
332 363
10 1 29 0 0 8320 0 19 15 0 0 4
272 395
324 395
324 326
332 326
1 6 30 0 0 8192 0 3 20 0 0 4
159 442
181 442
181 209
209 209
1 5 30 0 0 8320 0 3 20 0 0 4
159 442
181 442
181 200
209 200
1 8 30 0 0 0 0 3 20 0 0 4
159 442
181 442
181 227
209 227
1 9 30 0 0 0 0 3 20 0 0 4
159 442
181 442
181 245
209 245
1 6 30 0 0 0 0 3 19 0 0 4
159 442
185 442
185 413
208 413
1 5 30 0 0 0 0 3 19 0 0 4
159 442
190 442
190 404
208 404
1 8 30 0 0 0 0 3 19 0 0 4
159 442
195 442
195 431
208 431
1 9 30 0 0 0 0 3 19 0 0 4
159 442
200 442
200 449
208 449
1 7 31 0 0 8320 0 4 19 0 0 4
164 229
195 229
195 422
208 422
1 7 31 0 0 0 0 4 20 0 0 4
164 229
201 229
201 218
209 218
1 4 32 0 0 4224 0 17 19 0 0 3
165 335
165 395
208 395
2 3 33 0 0 4224 0 17 19 0 0 3
159 335
159 386
208 386
3 2 34 0 0 8320 0 17 19 0 0 3
153 335
153 377
208 377
4 1 35 0 0 8320 0 17 19 0 0 3
147 335
147 368
208 368
1 4 36 0 0 4224 0 18 20 0 0 3
163 105
163 191
209 191
2 3 37 0 0 4224 0 18 20 0 0 3
157 105
157 182
209 182
3 2 38 0 0 4224 0 18 20 0 0 3
151 105
151 173
209 173
4 1 39 0 0 8320 0 18 20 0 0 3
145 105
145 164
209 164
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
403 109 592 133
413 117 581 133
21 XS-2 SUBTRACTOR (1'S)
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
