CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
13
13 Logic Switch~
5 118 298 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43383.1 0
0
13 Logic Switch~
5 120 201 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
43383.1 0
0
13 Logic Switch~
5 121 111 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
43383.1 0
0
14 Logic Display~
6 745 490 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3421 0 0
2
43383.1 0
0
14 Logic Display~
6 744 403 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8157 0 0
2
43383.1 0
0
8 2-In OR~
219 615 513 0 3 22
0 5 4 2
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
5572 0 0
2
43383.1 0
0
8 2-In OR~
219 616 428 0 3 22
0 6 5 3
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
8901 0 0
2
43383.1 0
0
9 2-In AND~
219 406 382 0 3 22
0 7 8 4
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U2C
-12 -7 9 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
7361 0 0
2
43383.1 0
0
9 2-In AND~
219 358 383 0 3 22
0 9 7 5
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U2B
-12 -7 9 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
4747 0 0
2
43383.1 0
0
9 2-In AND~
219 306 382 0 3 22
0 10 9 6
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U2A
-12 -7 9 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
972 0 0
2
43383.1 0
0
9 Inverter~
13 208 329 0 2 22
0 7 11
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3472 0 0
2
43383.1 0
0
9 Inverter~
13 208 230 0 2 22
0 8 10
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
9998 0 0
2
43383.1 0
0
9 Inverter~
13 207 138 0 2 22
0 9 12
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3536 0 0
2
43383.1 0
0
24
3 1 2 0 0 8336 0 6 4 0 0 4
648 513
648 519
745 519
745 508
3 1 3 0 0 4224 0 7 5 0 0 3
649 428
744 428
744 421
2 0 4 0 0 4224 0 6 0 0 7 2
602 522
404 522
1 0 5 0 0 4096 0 6 0 0 8 2
602 504
356 504
2 0 5 0 0 4224 0 7 0 0 8 2
603 437
356 437
1 0 6 0 0 4224 0 7 0 0 9 2
603 419
304 419
3 0 4 0 0 0 0 8 0 0 0 2
404 405
404 581
3 0 5 0 0 0 0 9 0 0 0 2
356 406
356 581
3 0 6 0 0 0 0 10 0 0 0 2
304 405
304 581
1 0 7 0 0 4096 0 8 0 0 22 2
413 360
413 298
2 0 8 0 0 4096 0 8 0 0 23 2
395 360
395 201
1 0 9 0 0 4096 0 9 0 0 24 2
365 361
365 111
2 0 7 0 0 4096 0 9 0 0 22 2
347 361
347 298
1 0 10 0 0 4096 0 10 0 0 18 2
313 360
313 230
2 0 9 0 0 0 0 10 0 0 24 2
295 360
295 111
2 0 11 0 0 4224 0 11 0 0 0 2
229 329
655 329
1 1 7 0 0 0 0 1 11 0 0 4
130 298
185 298
185 329
193 329
2 0 10 0 0 4224 0 12 0 0 0 2
229 230
655 230
1 1 8 0 0 0 0 2 12 0 0 4
132 201
185 201
185 230
193 230
2 0 12 0 0 4224 0 13 0 0 0 2
228 138
654 138
1 1 9 0 0 0 0 3 13 0 0 4
133 111
184 111
184 138
192 138
1 0 7 0 0 4224 0 1 0 0 0 2
130 298
655 298
1 0 8 0 0 4224 0 2 0 0 0 2
132 201
655 201
1 0 9 0 0 4224 0 3 0 0 0 2
133 111
655 111
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
786 475 823 499
796 483 812 499
2 F2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
785 390 822 414
795 398 811 414
2 F1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
64 278 93 302
74 286 82 302
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
64 183 93 207
74 191 82 207
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
65 92 94 116
75 100 83 116
1 A
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
