CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
40 40 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 E:\CM60S\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
143654930 0
0
6 Title:
5 Name:
0
0
0
24
13 Logic Switch~
5 465 232 0 1 11
0 5
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
43331.8 0
0
13 Logic Switch~
5 93 409 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
43331.8 1
0
13 Logic Switch~
5 94 363 0 1 11
0 16
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
43331.8 2
0
13 Logic Switch~
5 94 320 0 1 11
0 9
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
43331.8 3
0
13 Logic Switch~
5 95 210 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8157 0 0
2
43331.8 4
0
13 Logic Switch~
5 97 163 0 1 11
0 14
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
43331.8 5
0
13 Logic Switch~
5 99 114 0 1 11
0 10
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
43331.8 6
0
14 Logic Display~
6 813 243 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7361 0 0
2
43331.8 7
0
14 Logic Display~
6 813 296 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4747 0 0
2
43331.8 8
0
9 2-In AND~
219 230 558 0 3 22
0 10 9 8
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
972 0 0
2
43331.8 9
0
14 Logic Display~
6 814 347 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3472 0 0
2
43331.8 10
0
9 2-In AND~
219 230 497 0 3 22
0 14 9 13
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
9998 0 0
2
43331.8 11
0
9 2-In AND~
219 229 445 0 3 22
0 10 16 15
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
3536 0 0
2
43331.8 12
0
14 Logic Display~
6 815 401 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4597 0 0
2
43331.8 13
0
9 2-In AND~
219 230 392 0 3 22
0 19 9 18
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3835 0 0
2
43331.8 14
0
6 74LS83
105 572 220 0 14 29
0 4 7 12 18 5 5 5 20 5
3 6 11 17 2
0
0 0 13024 0
7 74LS83A
-24 -60 25 -52
2 U4
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
3670 0 0
2
43331.8 15
0
9 2-In AND~
219 231 336 0 3 22
0 14 16 21
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
5616 0 0
2
43331.8 16
0
9 2-In AND~
219 231 283 0 3 22
0 10 23 22
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
9323 0 0
2
43331.8 17
0
14 Logic Display~
6 816 461 0 1 2
10 24
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
317 0 0
2
43331.8 18
0
9 2-In AND~
219 231 105 0 3 22
0 14 23 26
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3108 0 0
2
43331.8 19
0
9 2-In AND~
219 231 163 0 3 22
0 19 16 25
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
4299 0 0
2
43331.8 20
0
14 Logic Display~
6 816 521 0 1 2
10 27
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9672 0 0
2
43331.8 21
0
9 2-In AND~
219 231 228 0 3 22
0 19 23 27
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
7876 0 0
2
43331.8 22
0
6 74LS83
105 466 105 0 14 29
0 8 15 22 26 5 13 21 25 5
7 12 20 24 4
0
0 0 13024 0
7 74LS83A
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
6369 0 0
2
43331.8 23
0
43
0 14 2 0 0 4224 0 0 16 0 0 3
605 266
605 265
604 265
10 1 3 0 0 4224 0 16 8 0 0 5
604 211
800 211
800 269
813 269
813 261
14 1 4 0 0 4224 0 24 16 0 0 4
498 150
532 150
532 184
540 184
1 9 5 0 0 12288 0 1 24 0 0 6
477 232
502 232
502 165
426 165
426 150
434 150
1 9 5 0 0 0 0 1 16 0 0 4
477 232
532 232
532 265
540 265
1 5 5 0 0 0 0 1 16 0 0 4
477 232
532 232
532 220
540 220
11 1 6 0 0 4224 0 16 9 0 0 5
604 220
800 220
800 322
813 322
813 314
1 6 5 0 0 0 0 1 16 0 0 4
477 232
532 232
532 229
540 229
10 2 7 0 0 8320 0 24 16 0 0 4
498 96
532 96
532 193
540 193
1 5 5 0 0 8320 0 1 24 0 0 6
477 232
502 232
502 49
426 49
426 105
434 105
3 1 8 0 0 8320 0 10 24 0 0 4
251 558
426 558
426 69
434 69
1 2 9 0 0 8320 0 4 10 0 0 4
106 320
198 320
198 567
206 567
1 1 10 0 0 8320 0 7 10 0 0 4
111 114
198 114
198 549
206 549
12 1 11 0 0 4224 0 16 11 0 0 5
604 229
801 229
801 373
814 373
814 365
1 7 5 0 0 0 0 1 16 0 0 4
477 232
532 232
532 238
540 238
11 3 12 0 0 8320 0 24 16 0 0 4
498 105
532 105
532 202
540 202
3 6 13 0 0 8320 0 12 24 0 0 4
251 497
426 497
426 114
434 114
1 2 9 0 0 0 0 4 12 0 0 4
106 320
198 320
198 506
206 506
1 1 14 0 0 8320 0 6 12 0 0 4
109 163
198 163
198 488
206 488
3 2 15 0 0 8320 0 13 24 0 0 4
250 445
426 445
426 78
434 78
1 2 16 0 0 4096 0 3 13 0 0 4
106 363
197 363
197 454
205 454
1 1 10 0 0 0 0 7 13 0 0 4
111 114
197 114
197 436
205 436
13 1 17 0 0 4224 0 16 14 0 0 5
604 238
802 238
802 427
815 427
815 419
3 4 18 0 0 4224 0 15 16 0 0 4
251 392
532 392
532 211
540 211
1 2 9 0 0 0 0 4 15 0 0 4
106 320
198 320
198 401
206 401
1 1 19 0 0 8320 0 5 15 0 0 4
107 210
198 210
198 383
206 383
12 8 20 0 0 8320 0 24 16 0 0 4
498 114
532 114
532 247
540 247
3 7 21 0 0 8320 0 17 24 0 0 4
252 336
426 336
426 123
434 123
3 3 22 0 0 8320 0 18 24 0 0 4
252 283
426 283
426 87
434 87
1 2 16 0 0 4096 0 3 17 0 0 4
106 363
199 363
199 345
207 345
1 1 14 0 0 0 0 6 17 0 0 4
109 163
199 163
199 327
207 327
1 2 23 0 0 8192 0 2 18 0 0 4
105 409
199 409
199 292
207 292
1 1 10 0 0 0 0 7 18 0 0 4
111 114
199 114
199 274
207 274
13 1 24 0 0 8320 0 24 19 0 0 5
498 123
803 123
803 487
816 487
816 479
3 8 25 0 0 4224 0 21 24 0 0 4
252 163
426 163
426 132
434 132
3 4 26 0 0 4224 0 20 24 0 0 4
252 105
426 105
426 96
434 96
1 2 16 0 0 8320 0 3 21 0 0 4
106 363
199 363
199 172
207 172
1 1 19 0 0 0 0 5 21 0 0 4
107 210
199 210
199 154
207 154
1 2 23 0 0 8320 0 2 20 0 0 4
105 409
199 409
199 114
207 114
1 1 14 0 0 0 0 6 20 0 0 4
109 163
199 163
199 96
207 96
3 1 27 0 0 12416 0 23 22 0 0 5
252 228
433 228
433 547
816 547
816 539
1 2 23 0 0 0 0 2 23 0 0 4
105 409
199 409
199 237
207 237
1 1 19 0 0 0 0 5 23 0 0 4
107 210
199 210
199 219
207 219
13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
429 602 578 624
439 609 567 625
16 3 BIT MULTIPLIER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
52 93 76 117
62 101 78 117
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
49 142 73 166
59 150 75 166
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
46 190 70 214
56 198 72 214
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
44 290 68 314
54 298 70 314
2 B2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
45 337 69 361
55 345 71 361
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
43 385 67 409
53 393 69 409
2 B0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
821 509 845 533
831 517 847 533
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
821 449 845 473
831 457 847 473
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
820 392 844 416
830 400 846 416
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
816 336 840 360
826 344 842 360
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
817 287 841 311
827 295 843 311
2 S4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
816 233 840 257
826 241 842 257
2 S5
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
