CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
20 10 30 80 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
22
13 Logic Switch~
5 35 349 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43353.9 0
0
13 Logic Switch~
5 34 540 0 1 11
0 27
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
43353.9 0
0
13 Logic Switch~
5 35 585 0 1 11
0 29
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
43353.9 0
0
13 Logic Switch~
5 34 441 0 1 11
0 28
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3421 0 0
2
43353.9 0
0
13 Logic Switch~
5 32 489 0 1 11
0 30
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8157 0 0
2
43353.9 0
0
12 Hex Display~
7 127 682 0 16 19
10 9 8 7 6 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP5
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
5572 0 0
2
43354 0
0
12 Hex Display~
7 81 682 0 16 19
10 5 4 3 2 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP4
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
8901 0 0
2
43354 0
0
12 Hex Display~
7 614 48 0 18 19
10 15 16 17 18 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
7361 0 0
2
43354 0
0
12 Hex Display~
7 571 49 0 18 19
10 11 12 13 14 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
4747 0 0
2
43354 0
0
12 Hex Display~
7 530 49 0 16 19
10 10 63 64 65 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 0 0 0 0
4 DISP
972 0 0
2
43354 0
0
6 74LS93
109 131 577 0 8 17
0 27 27 29 5 2 3 4 5
0
0 0 4848 0
6 74LS93
-21 -35 21 -27
3 U10
-11 -36 10 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 0 0 0 0
1 U
3472 0 0
2
43353.9 0
0
6 74LS93
109 133 478 0 8 17
0 28 28 30 9 6 7 8 9
0
0 0 4848 0
6 74LS93
-21 -35 21 -27
2 U9
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 0 0 0 0
1 U
9998 0 0
2
43353.9 0
0
8 Hex Key~
166 252 52 0 11 12
0 35 36 37 38 0 0 0 0 0
1 49
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
3536 0 0
2
43353.9 0
0
8 Hex Key~
166 202 53 0 11 12
0 31 32 33 34 0 0 0 0 0
1 49
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
4597 0 0
2
43353.9 0
0
2 FA
94 386 102 0 5 11
0 38 6 24 20 18
2 FA
1 0 688 0
0
2 U1
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
3835 0 0
2
43334.9 0
0
2 FA
94 386 179 0 5 11
0 37 7 25 24 17
2 FA
2 0 688 0
0
2 U2
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
3670 0 0
2
43334.9 0
0
2 FA
94 386 256 0 5 11
0 36 8 26 25 16
2 FA
3 0 688 0
0
2 U3
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
5616 0 0
2
43334.9 0
0
2 FA
94 385 335 0 5 11
0 35 9 19 26 15
2 FA
4 0 688 0
0
2 U4
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
9323 0 0
2
43334.9 0
0
2 FA
94 384 415 0 5 11
0 34 2 23 10 14
2 FA
5 0 688 0
0
2 U5
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
317 0 0
2
43334.9 0
0
2 FA
94 384 498 0 5 11
0 33 3 22 23 13
2 FA
6 0 688 0
0
2 U6
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
3108 0 0
2
43334.9 0
0
2 FA
94 383 588 0 5 11
0 32 4 21 22 12
2 FA
7 0 688 0
0
2 U7
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
4299 0 0
2
43334.9 0
0
2 FA
94 383 675 0 5 11
0 31 5 20 21 11
2 FA
8 0 688 0
0
2 U8
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
9672 0 0
2
43334.9 0
0
49
5 4 2 0 0 8320 0 11 7 0 0 5
163 568
217 568
217 749
72 749
72 706
6 3 3 0 0 8192 0 11 7 0 0 5
163 577
202 577
202 744
78 744
78 706
7 2 4 0 0 8192 0 11 7 0 0 5
163 586
197 586
197 739
84 739
84 706
8 1 5 0 0 8192 0 11 7 0 0 5
163 595
167 595
167 734
90 734
90 706
5 4 6 0 0 8192 0 12 6 0 0 5
165 469
194 469
194 729
118 729
118 706
6 3 7 0 0 8192 0 12 6 0 0 5
165 478
189 478
189 724
124 724
124 706
7 2 8 0 0 8320 0 12 6 0 0 5
165 487
184 487
184 719
130 719
130 706
8 1 9 0 0 8320 0 12 6 0 0 5
165 496
179 496
179 714
136 714
136 706
4 1 10 0 0 8320 0 19 10 0 0 3
417 433
539 433
539 73
5 1 11 0 0 8320 0 22 9 0 0 3
416 675
580 675
580 73
5 2 12 0 0 8320 0 21 9 0 0 3
416 588
574 588
574 73
5 3 13 0 0 8320 0 20 9 0 0 3
417 498
568 498
568 73
5 4 14 0 0 8320 0 19 9 0 0 3
417 415
562 415
562 73
5 1 15 0 0 8320 0 18 8 0 0 3
418 335
623 335
623 72
5 2 16 0 0 4224 0 17 8 0 0 3
419 256
617 256
617 72
5 3 17 0 0 4224 0 16 8 0 0 3
419 179
611 179
611 72
5 4 18 0 0 4224 0 15 8 0 0 3
419 102
605 102
605 72
1 3 19 0 0 4224 0 1 18 0 0 4
47 349
324 349
324 353
352 353
4 3 20 0 0 8320 0 15 22 0 0 6
419 120
432 120
432 717
342 717
342 693
350 693
4 3 21 0 0 12416 0 22 21 0 0 5
416 693
421 693
421 635
350 635
350 606
4 3 22 0 0 12416 0 21 20 0 0 6
416 606
421 606
421 530
338 530
338 516
351 516
4 3 23 0 0 12416 0 20 19 0 0 5
417 516
423 516
423 458
351 458
351 433
4 3 24 0 0 12416 0 16 15 0 0 6
419 197
423 197
423 140
345 140
345 120
353 120
4 3 25 0 0 12416 0 17 16 0 0 6
419 274
423 274
423 218
345 218
345 197
353 197
4 3 26 0 0 12416 0 18 17 0 0 6
418 353
423 353
423 288
345 288
345 274
353 274
5 2 2 0 0 128 0 11 19 0 0 4
163 568
323 568
323 424
351 424
6 2 3 0 0 4224 0 11 20 0 0 4
163 577
343 577
343 507
351 507
7 2 4 0 0 4224 0 11 21 0 0 4
163 586
337 586
337 597
350 597
8 2 5 0 0 4224 0 11 22 0 0 4
163 595
342 595
342 684
350 684
5 2 6 0 0 8320 0 12 15 0 0 4
165 469
330 469
330 111
353 111
6 2 7 0 0 8320 0 12 16 0 0 4
165 478
335 478
335 188
353 188
7 2 8 0 0 128 0 12 17 0 0 4
165 487
340 487
340 265
353 265
8 2 9 0 0 144 0 12 18 0 0 5
165 496
165 494
344 494
344 344
352 344
4 8 5 0 0 0 0 11 11 0 0 6
93 595
89 595
89 610
171 610
171 595
163 595
4 8 9 0 0 0 0 12 12 0 0 6
95 496
91 496
91 511
173 511
173 496
165 496
1 2 27 0 0 8192 0 2 11 0 0 4
46 540
80 540
80 577
99 577
1 1 27 0 0 4224 0 2 11 0 0 4
46 540
85 540
85 568
99 568
1 2 28 0 0 8192 0 4 12 0 0 4
46 441
82 441
82 478
101 478
1 1 28 0 0 4224 0 4 12 0 0 4
46 441
87 441
87 469
101 469
1 3 29 0 0 4224 0 3 11 0 0 4
47 585
85 585
85 586
93 586
1 3 30 0 0 4224 0 5 12 0 0 4
44 489
87 489
87 487
95 487
1 1 31 0 0 4224 0 14 22 0 0 3
211 77
211 675
350 675
2 1 32 0 0 4224 0 14 21 0 0 3
205 77
205 588
350 588
3 1 33 0 0 4224 0 14 20 0 0 3
199 77
199 498
351 498
4 1 34 0 0 4224 0 14 19 0 0 3
193 77
193 415
351 415
1 1 35 0 0 4224 0 13 18 0 0 3
261 76
261 335
352 335
2 1 36 0 0 4224 0 13 17 0 0 3
255 76
255 256
353 256
3 1 37 0 0 8320 0 13 16 0 0 3
249 76
249 179
353 179
4 1 38 0 0 8320 0 13 15 0 0 3
243 76
243 102
353 102
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
