CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
10 10 30 60 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
28
13 Logic Switch~
5 63 486 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43335.1 0
0
13 Logic Switch~
5 63 353 0 10 11
0 29 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 64 294 0 10 11
0 27 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3124 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 66 239 0 10 11
0 25 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 67 151 0 10 11
0 28 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8157 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 69 96 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5572 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 70 45 0 10 11
0 24 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8901 0 0
2
5.89859e-315 0
0
14 Logic Display~
6 954 842 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7361 0 0
2
43335.1 0
0
14 Logic Display~
6 864 844 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4747 0 0
2
43335.1 0
0
14 Logic Display~
6 675 847 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
972 0 0
2
43335.1 0
0
14 Logic Display~
6 457 849 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3472 0 0
2
43335.1 0
0
14 Logic Display~
6 300 851 0 1 2
10 20
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9998 0 0
2
43335.1 0
0
14 Logic Display~
6 158 855 0 1 2
10 23
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3536 0 0
2
43335.1 0
0
9 2-In AND~
219 789 394 0 3 22
0 24 25 6
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U11A
-15 -11 13 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
4597 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 587 394 0 3 22
0 25 26 12
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3D
-12 -11 9 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
3835 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 549 395 0 3 22
0 27 24 13
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3C
-12 -11 9 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
3670 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 398 396 0 3 22
0 25 28 19
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3B
-12 -11 9 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
5616 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 358 396 0 3 22
0 27 26 18
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3A
-12 -11 9 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
9323 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 317 397 0 3 22
0 29 24 17
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1D
-12 -11 9 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
317 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 213 396 0 3 22
0 27 28 22
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1C
-12 -11 9 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3108 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 169 396 0 3 22
0 29 26 21
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1B
-12 -10 9 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
4299 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 121 397 0 3 22
0 28 29 23
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1A
-12 -10 9 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
9672 0 0
2
5.89859e-315 0
0
2 FA
94 190 472 0 5 11
0 22 21 8 15 20
2 FA
10 0 688 0
0
2 U2
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
7876 0 0
2
43334.9 0
0
2 FA
94 359 470 0 5 11
0 19 18 17 11 16
2 FA
11 0 688 0
0
2 U4
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
6369 0 0
2
43334.9 0
0
2 FA
94 359 568 0 5 11
0 15 16 8 9 14
2 FA
12 0 688 0
0
2 U5
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
9172 0 0
2
43334.9 0
0
2 FA
94 569 470 0 5 11
0 12 13 11 5 10
2 FA
13 0 688 0
0
2 U6
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
7100 0 0
2
43334.9 0
0
2 FA
94 570 568 0 5 11
0 9 10 8 4 7
2 FA
14 0 688 0
0
2 U7
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
3820 0 0
2
43334.9 0
0
2 FA
94 788 469 0 5 11
0 6 4 5 2 3
2 FA
15 0 688 0
0
2 U8
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
7678 0 0
2
43334.9 0
0
48
4 1 2 0 0 8320 0 28 8 0 0 5
821 487
930 487
930 889
954 889
954 860
5 1 3 0 0 8320 0 28 9 0 0 5
821 469
839 469
839 889
864 889
864 862
4 2 4 0 0 4224 0 27 28 0 0 4
603 586
722 586
722 478
755 478
4 3 5 0 0 8320 0 26 28 0 0 3
602 488
602 487
755 487
3 1 6 0 0 8320 0 14 28 0 0 5
787 417
787 428
732 428
732 469
755 469
5 1 7 0 0 8320 0 27 10 0 0 5
603 568
641 568
641 889
675 889
675 865
0 3 8 0 0 8320 0 0 27 14 0 7
159 586
159 608
463 608
463 593
528 593
528 586
537 586
4 1 9 0 0 4224 0 25 27 0 0 4
392 586
515 586
515 568
537 568
5 2 10 0 0 12416 0 26 27 0 0 6
602 470
642 470
642 521
489 521
489 577
537 577
4 3 11 0 0 4224 0 24 26 0 0 2
392 488
536 488
3 1 12 0 0 8320 0 15 26 0 0 5
585 417
585 430
505 430
505 470
536 470
3 2 13 0 0 8320 0 16 26 0 0 4
547 418
494 418
494 479
536 479
5 1 14 0 0 8320 0 25 11 0 0 5
392 568
419 568
419 889
457 889
457 867
1 3 8 0 0 0 0 1 25 0 0 3
75 486
75 586
326 586
4 1 15 0 0 8320 0 23 25 0 0 4
223 490
279 490
279 568
326 568
5 2 16 0 0 12416 0 24 25 0 0 6
392 470
419 470
419 522
291 522
291 577
326 577
3 3 17 0 0 4224 0 19 24 0 0 3
315 420
315 488
326 488
3 2 18 0 0 8320 0 18 24 0 0 5
356 419
356 430
290 430
290 479
326 479
3 1 19 0 0 8320 0 17 24 0 0 5
396 419
396 437
299 437
299 470
326 470
5 1 20 0 0 8320 0 23 12 0 0 5
223 472
251 472
251 889
300 889
300 869
1 3 8 0 0 16 0 1 23 0 0 3
75 486
75 490
157 490
3 2 21 0 0 12416 0 21 23 0 0 5
167 419
167 431
136 431
136 481
157 481
3 1 22 0 0 8320 0 20 23 0 0 5
211 419
211 437
143 437
143 472
157 472
3 1 23 0 0 4224 0 22 13 0 0 4
119 420
119 889
158 889
158 873
1 0 24 0 0 4096 0 14 0 0 48 2
796 372
796 45
2 0 25 0 0 4096 0 14 0 0 45 2
778 372
778 239
1 0 25 0 0 0 0 15 0 0 45 2
594 372
594 239
2 0 26 0 0 4096 0 15 0 0 47 2
576 372
576 96
1 0 27 0 0 4096 0 16 0 0 44 2
556 373
556 294
2 0 24 0 0 4096 0 16 0 0 48 2
538 373
538 45
1 0 25 0 0 4096 0 17 0 0 45 2
405 374
405 239
2 0 28 0 0 4096 0 17 0 0 46 2
387 374
387 151
1 0 27 0 0 4096 0 18 0 0 44 2
365 374
365 294
2 0 26 0 0 4096 0 18 0 0 47 2
347 374
347 96
1 0 29 0 0 4096 0 19 0 0 43 2
324 375
324 353
2 0 24 0 0 4096 0 19 0 0 48 2
306 375
306 45
1 0 27 0 0 0 0 20 0 0 44 2
220 374
220 294
2 0 28 0 0 0 0 20 0 0 46 2
202 374
202 151
1 0 29 0 0 0 0 21 0 0 43 2
176 374
176 353
2 0 26 0 0 0 0 21 0 0 47 2
158 374
158 96
1 0 28 0 0 4096 0 22 0 0 46 2
128 375
128 151
2 0 29 0 0 0 0 22 0 0 43 2
110 375
110 353
1 0 29 0 0 4224 0 2 0 0 0 2
75 353
1156 353
1 0 27 0 0 4224 0 3 0 0 0 2
76 294
1155 294
1 0 25 0 0 4224 0 4 0 0 0 2
78 239
1156 239
1 0 28 0 0 4224 0 5 0 0 0 2
79 151
1156 151
1 0 26 0 0 4224 0 6 0 0 0 2
81 96
1155 96
1 0 24 0 0 4224 0 7 0 0 0 2
82 45
1155 45
12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
936 775 973 799
946 783 962 799
2 S5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
846 782 883 806
856 790 872 806
2 S4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
656 785 693 809
666 793 682 809
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
439 781 476 805
449 789 465 805
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
282 782 319 806
292 790 308 806
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
140 786 177 810
150 794 166 810
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
20 23 57 47
30 31 46 47
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
20 74 57 98
30 82 46 98
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
19 127 56 151
29 135 45 151
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
18 215 55 239
28 223 44 239
2 B2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
17 273 54 297
27 281 43 297
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
16 329 53 353
26 337 42 353
2 B0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
