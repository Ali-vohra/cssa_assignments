CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
15
13 Logic Switch~
5 541 560 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V3
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3670 0 0
2
5.89862e-315 0
0
13 Logic Switch~
5 608 559 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V4
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5616 0 0
2
5.89862e-315 0
0
13 Logic Switch~
5 456 560 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V2
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9323 0 0
2
5.89862e-315 5.30499e-315
0
13 Logic Switch~
5 128 255 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
317 0 0
2
5.89862e-315 5.32571e-315
0
9 Inverter~
13 423 506 0 2 22
0 8 9
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U3A
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3108 0 0
2
5.89862e-315 5.34643e-315
0
14 Logic Display~
6 706 394 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4299 0 0
2
5.89862e-315 5.3568e-315
0
14 Logic Display~
6 706 343 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9672 0 0
2
5.89862e-315 5.36716e-315
0
14 Logic Display~
6 706 291 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7876 0 0
2
5.89862e-315 5.37752e-315
0
14 Logic Display~
6 703 237 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6369 0 0
2
5.89862e-315 5.38788e-315
0
14 Logic Display~
6 702 186 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9172 0 0
2
5.89862e-315 5.39306e-315
0
14 Logic Display~
6 703 134 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7100 0 0
2
5.89862e-315 5.39824e-315
0
14 Logic Display~
6 702 84 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3820 0 0
2
5.89862e-315 5.40342e-315
0
14 Logic Display~
6 702 36 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7678 0 0
2
5.89862e-315 5.4086e-315
0
10 4x1 DEMUX~
94 341 136 0 8 17
0 14 13 12 11 10 2 7 8
10 4x1 DEMUX~
3 0 560 0
0
2 U1
1 -68 15 -60
0
0
0
0
0
0
17

0 4 9 10 11 12 14 15 16 4
9 10 11 12 14 15 16 0
0 0 0 0 0 0 0 0
1 U
961 0 0
2
43362 0
0
10 4x1 DEMUX~
94 342 344 0 8 17
0 14 3 4 5 6 2 7 9
10 4x1 DEMUX~
4 0 560 0
0
2 U2
1 -68 15 -60
0
0
0
0
0
0
17

0 4 9 10 11 12 14 15 16 4
9 10 11 12 14 15 16 0
0 0 0 0 0 0 0 0
1 U
3178 0 0
2
43362 0
0
17
1 6 2 0 0 4224 0 1 14 0 0 3
542 547
542 125
390 125
1 6 2 0 0 0 0 1 15 0 0 3
542 547
542 333
391 333
2 1 3 0 0 4224 0 15 9 0 0 5
391 390
684 390
684 263
703 263
703 255
3 1 4 0 0 4224 0 15 8 0 0 5
391 379
688 379
688 317
706 317
706 309
4 1 5 0 0 4224 0 15 7 0 0 3
391 367
706 367
706 361
5 1 6 0 0 4224 0 15 6 0 0 5
391 355
694 355
694 420
706 420
706 412
1 7 7 0 0 4096 0 2 15 0 0 3
609 546
609 321
391 321
1 7 7 0 0 4224 0 2 14 0 0 3
609 546
609 113
390 113
1 8 8 0 0 4224 0 3 14 0 0 3
457 547
457 101
390 101
2 8 9 0 0 4224 0 5 15 0 0 3
426 488
426 309
391 309
1 1 8 0 0 0 0 3 5 0 0 4
457 547
457 532
426 532
426 524
5 1 10 0 0 4224 0 14 10 0 0 5
390 147
679 147
679 212
702 212
702 204
4 1 11 0 0 4224 0 14 11 0 0 3
390 159
703 159
703 152
3 1 12 0 0 4224 0 14 12 0 0 5
390 171
685 171
685 110
702 110
702 102
2 1 13 0 0 4224 0 14 13 0 0 5
390 182
690 182
690 62
702 62
702 54
1 1 14 0 0 4096 0 15 4 0 0 4
309 344
154 344
154 255
140 255
1 1 14 0 0 4224 0 14 4 0 0 4
308 136
149 136
149 255
140 255
12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
525 576 562 600
535 584 551 600
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
65 232 102 256
75 240 91 256
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
440 581 477 605
450 589 466 605
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
594 579 631 603
604 587 620 603
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
726 21 763 45
736 29 752 45
2 D7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
725 70 762 94
735 78 751 94
2 D6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
726 120 763 144
736 128 752 144
2 D5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
724 172 761 196
734 180 750 196
2 D4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
723 222 760 246
733 230 749 246
2 D3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
724 275 761 299
734 283 750 299
2 D2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
726 328 763 352
736 336 752 352
2 D1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
722 378 759 402
732 386 748 402
2 D0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
