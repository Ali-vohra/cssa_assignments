CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
340 100 3 160 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
10
12 Hex Display~
7 604 58 0 18 19
10 2 3 4 5 0 0 0 0 0
0 1 0 1 1 0 1 1 5
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
5130 0 0
2
5.89855e-315 0
0
12 Hex Display~
7 384 63 0 16 19
10 6 7 8 9 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
391 0 0
2
5.89855e-315 0
0
5 4071~
219 509 201 0 3 22
0 11 12 10
0
0 0 608 180
4 4071
-7 -24 21 -16
3 U4A
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
3124 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 399 148 0 3 22
0 13 14 12
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U3D
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
3421 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 607 153 0 3 22
0 4 3 14
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U3C
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
8157 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 398 217 0 3 22
0 8 8 13
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U3B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
5572 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 606 209 0 3 22
0 5 3 11
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U3A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
8901 0 0
2
5.89855e-315 0
0
7 Pulser~
4 516 367 0 10 12
0 16 17 15 18 0 0 5 5 2
7
0
0 0 4640 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7361 0 0
2
5.89855e-315 0
0
6 74LS93
109 599 285 0 8 17
0 10 10 15 2 5 4 3 2
0
0 0 4832 0
6 74LS93
-21 -35 21 -27
2 U2
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
4747 0 0
2
5.89855e-315 0
0
6 74LS93
109 393 287 0 8 17
0 12 12 5 6 9 8 7 6
0
0 0 4832 0
6 74LS93
-21 -35 21 -27
2 U1
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
972 0 0
2
5.89855e-315 0
0
26
8 1 2 0 0 8320 0 9 1 0 0 5
631 303
675 303
675 105
613 105
613 82
7 2 3 0 0 8320 0 9 1 0 0 5
631 294
670 294
670 100
607 100
607 82
6 3 4 0 0 8320 0 9 1 0 0 5
631 285
665 285
665 95
601 95
601 82
5 4 5 0 0 8192 0 9 1 0 0 5
631 276
660 276
660 90
595 90
595 82
8 1 6 0 0 8320 0 10 2 0 0 5
425 305
454 305
454 110
393 110
393 87
7 2 7 0 0 8320 0 10 2 0 0 5
425 296
449 296
449 105
387 105
387 87
6 3 8 0 0 8320 0 10 2 0 0 5
425 287
444 287
444 100
381 100
381 87
5 4 9 0 0 8320 0 10 2 0 0 5
425 278
439 278
439 95
375 95
375 87
0 2 10 0 0 8192 0 0 9 10 0 3
513 276
513 285
567 285
3 1 10 0 0 8320 0 3 9 0 0 3
482 201
482 276
567 276
1 3 11 0 0 8320 0 3 7 0 0 3
528 210
528 209
579 209
3 2 12 0 0 8320 0 4 3 0 0 5
372 148
372 118
539 118
539 192
528 192
3 2 12 0 0 0 0 4 10 0 0 4
372 148
342 148
342 287
361 287
3 1 12 0 0 0 0 4 10 0 0 4
372 148
347 148
347 278
361 278
3 1 13 0 0 8320 0 6 4 0 0 6
371 217
370 217
370 128
432 128
432 157
417 157
3 2 14 0 0 4224 0 5 4 0 0 4
580 153
427 153
427 139
417 139
7 2 3 0 0 0 0 9 5 0 0 4
631 294
655 294
655 144
625 144
6 1 4 0 0 0 0 9 5 0 0 4
631 285
650 285
650 162
625 162
6 2 8 0 0 0 0 10 6 0 0 4
425 287
434 287
434 208
416 208
6 1 8 0 0 0 0 10 6 0 0 4
425 287
429 287
429 226
416 226
7 2 3 0 0 0 0 9 7 0 0 4
631 294
646 294
646 200
624 200
5 1 5 0 0 0 0 9 7 0 0 4
631 276
636 276
636 218
624 218
8 4 6 0 0 0 0 10 10 0 0 6
425 305
429 305
429 320
342 320
342 305
355 305
5 3 5 0 0 12416 0 9 10 0 0 6
631 276
640 276
640 325
347 325
347 296
355 296
8 4 2 0 0 0 0 9 9 0 0 6
631 303
635 303
635 318
548 318
548 303
561 303
3 3 15 0 0 8320 0 8 9 0 0 4
540 358
553 358
553 294
561 294
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
418 397 591 421
424 402 584 418
20 DIVIDE BY 45 COUNTER
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
