CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
160 70 30 110 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 307 331 0 1 11
0 7
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 204 610 0 1 11
0 8
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89855e-315 0
0
14 Logic Display~
6 782 319 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3124 0 0
2
5.89855e-315 0
0
12 Hex Display~
7 678 183 0 18 19
10 3 4 5 6 0 0 0 0 0
0 1 1 1 1 1 1 1 8
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3421 0 0
2
5.89855e-315 0
0
5 4030~
219 243 520 0 3 22
0 13 8 9
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U2D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 1 0
1 U
8157 0 0
2
5.89855e-315 0
0
5 4030~
219 243 467 0 3 22
0 14 8 10
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U2C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 1 0
1 U
5572 0 0
2
5.89855e-315 0
0
5 4030~
219 243 416 0 3 22
0 15 8 11
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U2B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
8901 0 0
2
5.89855e-315 0
0
5 4030~
219 243 363 0 3 22
0 16 8 12
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U2A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
7361 0 0
2
5.89855e-315 0
0
8 Hex Key~
166 182 181 0 11 12
0 13 14 15 16 0 0 0 0 0
2 50
0
0 0 4640 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
4747 0 0
2
5.89855e-315 0
0
8 Hex Key~
166 288 183 0 11 12
0 17 18 19 20 0 0 0 0 0
6 54
0
0 0 4640 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
972 0 0
2
5.89855e-315 0
0
6 74LS83
105 423 288 0 14 29
0 20 19 18 17 12 11 10 9 7
6 5 4 3 2
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
3472 0 0
2
5.89855e-315 0
0
22
14 1 2 0 0 4224 0 11 3 0 0 5
455 333
770 333
770 345
782 345
782 337
13 1 3 0 0 4224 0 11 4 0 0 3
455 306
687 306
687 207
12 2 4 0 0 4224 0 11 4 0 0 3
455 297
681 297
681 207
11 3 5 0 0 4224 0 11 4 0 0 3
455 288
675 288
675 207
10 4 6 0 0 4224 0 11 4 0 0 3
455 279
669 279
669 207
1 9 7 0 0 4224 0 1 11 0 0 4
319 331
363 331
363 333
391 333
1 2 8 0 0 8320 0 2 8 0 0 4
216 610
221 610
221 372
227 372
1 2 8 0 0 0 0 2 7 0 0 4
216 610
221 610
221 425
227 425
1 2 8 0 0 0 0 2 6 0 0 4
216 610
221 610
221 476
227 476
1 2 8 0 0 0 0 2 5 0 0 4
216 610
221 610
221 529
227 529
3 8 9 0 0 8320 0 5 11 0 0 4
276 520
368 520
368 315
391 315
3 7 10 0 0 8320 0 6 11 0 0 4
276 467
373 467
373 306
391 306
3 6 11 0 0 8320 0 7 11 0 0 4
276 416
378 416
378 297
391 297
3 5 12 0 0 4224 0 8 11 0 0 4
276 363
383 363
383 288
391 288
1 1 13 0 0 4224 0 9 5 0 0 3
191 205
191 511
227 511
2 1 14 0 0 4224 0 9 6 0 0 3
185 205
185 458
227 458
3 1 15 0 0 4224 0 9 7 0 0 3
179 205
179 407
227 407
4 1 16 0 0 4224 0 9 8 0 0 3
173 205
173 354
227 354
1 4 17 0 0 8320 0 10 11 0 0 3
297 207
297 279
391 279
2 3 18 0 0 8320 0 10 11 0 0 3
291 207
291 270
391 270
3 2 19 0 0 8320 0 10 11 0 0 3
285 207
285 261
391 261
4 1 20 0 0 8320 0 10 11 0 0 3
279 207
279 252
391 252
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
373 78 518 99
381 84 509 99
16 BINARY ADDER/SUB
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
