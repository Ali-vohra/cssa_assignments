CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
40
13 Logic Switch~
5 189 820 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43354 0
0
13 Logic Switch~
5 139 821 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
391 0 0
2
43354 0
0
13 Logic Switch~
5 35 349 0 1 11
0 43
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89861e-315 0
0
13 Logic Switch~
5 34 540 0 1 11
0 51
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.89861e-315 0
0
13 Logic Switch~
5 35 585 0 1 11
0 53
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.89861e-315 0
0
13 Logic Switch~
5 34 441 0 1 11
0 52
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
5.89861e-315 0
0
13 Logic Switch~
5 32 489 0 1 11
0 54
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
5.89861e-315 0
0
9 Inverter~
13 325 1346 0 2 22
0 18 26
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U20B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
7361 0 0
2
43354 0
0
9 Inverter~
13 327 1260 0 2 22
0 19 27
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U20A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
4747 0 0
2
43354 0
0
9 Inverter~
13 327 1175 0 2 22
0 20 28
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U19F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
972 0 0
2
43354 0
0
9 Inverter~
13 327 1095 0 2 22
0 21 29
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U19E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
3472 0 0
2
43354 0
0
9 Inverter~
13 329 1012 0 2 22
0 22 30
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U19D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
9998 0 0
2
43354 0
0
9 Inverter~
13 329 930 0 2 22
0 23 31
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U19C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3536 0 0
2
43354 0
0
9 Inverter~
13 330 850 0 2 22
0 24 32
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U19B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
4597 0 0
2
43354 0
0
9 Inverter~
13 330 771 0 2 22
0 25 33
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U19A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3835 0 0
2
43354 0
0
12 Hex Display~
7 127 682 0 18 19
10 22 23 24 25 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP5
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3670 0 0
2
5.89861e-315 0
0
12 Hex Display~
7 81 682 0 18 19
10 18 19 20 21 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP4
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
5616 0 0
2
5.89861e-315 0
0
12 Hex Display~
7 614 48 0 16 19
10 39 40 41 42 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
9323 0 0
2
5.89861e-315 0
0
12 Hex Display~
7 571 49 0 18 19
10 35 36 37 38 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
317 0 0
2
5.89861e-315 0
0
12 Hex Display~
7 530 49 0 18 19
10 34 113 114 115 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
3108 0 0
2
5.89861e-315 0
0
6 74LS93
109 131 577 0 8 17
0 51 51 53 18 21 20 19 18
0
0 0 4848 0
6 74LS93
-21 -35 21 -27
3 U10
-11 -36 10 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
4299 0 0
2
5.89861e-315 0
0
6 74LS93
109 133 478 0 8 17
0 52 52 54 22 25 24 23 22
0
0 0 4848 0
6 74LS93
-21 -35 21 -27
2 U9
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
9672 0 0
2
5.89861e-315 0
0
8 Hex Key~
166 252 52 0 11 12
0 59 60 61 62 0 0 0 0 0
1 49
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
7876 0 0
2
5.89861e-315 0
0
8 Hex Key~
166 202 53 0 11 12
0 55 56 57 58 0 0 0 0 0
1 49
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
6369 0 0
2
5.89861e-315 0
0
2 FA
94 386 102 0 5 11
0 62 9 48 44 42
2 FA
1 0 688 0
0
2 U1
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 1 0 0 0
1 U
9172 0 0
2
5.89859e-315 0
0
2 FA
94 386 179 0 5 11
0 61 8 49 48 41
2 FA
2 0 688 0
0
2 U2
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 1 0 0 0
1 U
7100 0 0
2
5.89859e-315 0
0
2 FA
94 386 256 0 5 11
0 60 7 50 49 40
2 FA
3 0 688 0
0
2 U3
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 1 0 0 0
1 U
3820 0 0
2
5.89859e-315 0
0
2 FA
94 385 335 0 5 11
0 59 6 43 50 39
2 FA
4 0 688 0
0
2 U4
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 1 0 0 0
1 U
7678 0 0
2
5.89859e-315 0
0
2 FA
94 384 415 0 5 11
0 58 5 47 34 38
2 FA
5 0 688 0
0
2 U5
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 1 0 0 0
1 U
961 0 0
2
5.89859e-315 0
0
2 FA
94 384 498 0 5 11
0 57 4 46 47 37
2 FA
6 0 688 0
0
2 U6
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 1 0 0 0
1 U
3178 0 0
2
5.89859e-315 0
0
2 FA
94 383 588 0 5 11
0 56 3 45 46 36
2 FA
7 0 688 0
0
2 U7
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 1 0 0 0
1 U
3409 0 0
2
5.89859e-315 0
0
2 FA
94 383 675 0 5 11
0 55 2 44 45 35
2 FA
8 0 688 0
0
2 U8
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 1 0 0 0
1 U
3951 0 0
2
5.89859e-315 0
0
2 FA
94 384 771 0 5 11
0 33 13 14 87 9
2 FA
9 0 688 0
0
3 U11
-11 -29 10 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
8885 0 0
2
43334.9 0
0
2 FA
94 384 850 0 5 11
0 32 13 15 14 8
2 FA
10 0 688 0
0
3 U12
-11 -29 10 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
3780 0 0
2
43334.9 0
0
2 FA
94 384 930 0 5 11
0 31 13 16 15 7
2 FA
11 0 688 0
0
3 U13
-11 -29 10 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
9265 0 0
2
43334.9 0
0
2 FA
94 384 1012 0 5 11
0 30 17 13 16 6
2 FA
12 0 688 0
0
3 U14
-11 -29 10 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
9442 0 0
2
43334.9 0
0
2 FA
94 382 1095 0 5 11
0 29 13 10 100 5
2 FA
13 0 688 0
0
3 U15
-11 -29 10 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
9424 0 0
2
43334.9 0
0
2 FA
94 381 1175 0 5 11
0 28 13 11 10 4
2 FA
14 0 688 0
0
3 U16
-11 -29 10 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
9968 0 0
2
43334.9 0
0
2 FA
94 381 1260 0 5 11
0 27 13 12 11 3
2 FA
15 0 688 0
0
3 U17
-11 -29 10 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
9281 0 0
2
43334.9 0
0
2 FA
94 380 1346 0 5 11
0 26 17 13 12 2
2 FA
16 0 688 0
0
3 U18
-11 -29 10 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
8464 0 0
2
43334.9 0
0
81
5 2 2 0 0 8320 0 40 32 0 0 6
413 1346
511 1346
511 711
334 711
334 684
350 684
5 2 3 0 0 8320 0 39 31 0 0 6
414 1260
501 1260
501 628
341 628
341 597
350 597
5 2 4 0 0 8320 0 38 30 0 0 6
414 1175
491 1175
491 538
330 538
330 507
351 507
5 2 5 0 0 8320 0 37 29 0 0 6
415 1095
482 1095
482 452
345 452
345 424
351 424
5 2 6 0 0 8320 0 36 28 0 0 6
417 1012
472 1012
472 377
335 377
335 344
352 344
5 2 7 0 0 8320 0 35 27 0 0 6
417 930
461 930
461 296
335 296
335 265
353 265
5 2 8 0 0 8320 0 34 26 0 0 6
417 850
452 850
452 213
335 213
335 188
353 188
5 2 9 0 0 8320 0 33 25 0 0 6
417 771
442 771
442 146
341 146
341 111
353 111
4 3 10 0 0 12416 0 38 37 0 0 6
414 1193
433 1193
433 1135
340 1135
340 1113
349 1113
4 3 11 0 0 12416 0 39 38 0 0 6
414 1278
432 1278
432 1218
340 1218
340 1193
348 1193
4 3 12 0 0 12416 0 40 39 0 0 6
413 1364
431 1364
431 1304
339 1304
339 1278
348 1278
3 0 13 0 0 4096 0 36 0 0 19 2
351 1030
201 1030
0 3 13 0 0 0 0 0 40 17 0 3
201 1269
201 1364
347 1364
4 3 14 0 0 12416 0 34 33 0 0 6
417 868
433 868
433 810
343 810
343 789
351 789
4 3 15 0 0 12416 0 35 34 0 0 6
417 948
432 948
432 893
343 893
343 868
351 868
4 3 16 0 0 12416 0 36 35 0 0 6
417 1030
431 1030
431 972
344 972
344 948
351 948
0 2 13 0 0 0 0 0 39 18 0 3
201 1183
201 1269
348 1269
0 2 13 0 0 0 0 0 38 19 0 3
201 1104
201 1184
348 1184
1 2 13 0 0 4224 0 1 37 0 0 3
201 820
201 1104
349 1104
1 2 13 0 0 0 0 1 35 0 0 3
201 820
201 939
351 939
1 2 13 0 0 0 0 1 34 0 0 3
201 820
201 859
351 859
1 2 13 0 0 0 0 1 33 0 0 3
201 820
201 780
351 780
1 2 17 0 0 4224 0 2 40 0 0 3
151 821
151 1355
347 1355
1 2 17 0 0 0 0 2 36 0 0 3
151 821
151 1021
351 1021
8 1 18 0 0 8320 0 21 8 0 0 4
163 595
287 595
287 1346
310 1346
7 1 19 0 0 8320 0 21 9 0 0 4
163 586
279 586
279 1260
312 1260
6 1 20 0 0 8320 0 21 10 0 0 4
163 577
284 577
284 1175
312 1175
5 1 21 0 0 8320 0 21 11 0 0 4
163 568
299 568
299 1095
312 1095
8 1 22 0 0 8320 0 22 12 0 0 4
165 496
291 496
291 1012
314 1012
7 1 23 0 0 8320 0 22 13 0 0 4
165 487
296 487
296 930
314 930
6 1 24 0 0 8320 0 22 14 0 0 4
165 478
302 478
302 850
315 850
5 1 25 0 0 8320 0 22 15 0 0 4
165 469
307 469
307 771
315 771
2 1 26 0 0 8320 0 8 40 0 0 3
346 1346
346 1346
347 1346
2 1 27 0 0 0 0 9 39 0 0 2
348 1260
348 1260
2 1 28 0 0 0 0 10 38 0 0 2
348 1175
348 1175
2 1 29 0 0 4224 0 11 37 0 0 2
348 1095
349 1095
2 1 30 0 0 4224 0 12 36 0 0 2
350 1012
351 1012
2 1 31 0 0 4224 0 13 35 0 0 2
350 930
351 930
2 1 32 0 0 0 0 14 34 0 0 2
351 850
351 850
2 1 33 0 0 0 0 15 33 0 0 2
351 771
351 771
5 4 21 0 0 128 0 21 17 0 0 5
163 568
217 568
217 749
72 749
72 706
6 3 20 0 0 0 0 21 17 0 0 5
163 577
202 577
202 744
78 744
78 706
7 2 19 0 0 0 0 21 17 0 0 5
163 586
197 586
197 739
84 739
84 706
8 1 18 0 0 0 0 21 17 0 0 5
163 595
167 595
167 734
90 734
90 706
5 4 25 0 0 0 0 22 16 0 0 5
165 469
194 469
194 729
118 729
118 706
6 3 24 0 0 0 0 22 16 0 0 5
165 478
189 478
189 724
124 724
124 706
7 2 23 0 0 128 0 22 16 0 0 5
165 487
184 487
184 719
130 719
130 706
8 1 22 0 0 128 0 22 16 0 0 5
165 496
179 496
179 714
136 714
136 706
4 1 34 0 0 8320 0 29 20 0 0 3
417 433
539 433
539 73
5 1 35 0 0 8320 0 32 19 0 0 3
416 675
580 675
580 73
5 2 36 0 0 8320 0 31 19 0 0 3
416 588
574 588
574 73
5 3 37 0 0 8320 0 30 19 0 0 3
417 498
568 498
568 73
5 4 38 0 0 8320 0 29 19 0 0 3
417 415
562 415
562 73
5 1 39 0 0 8320 0 28 18 0 0 3
418 335
623 335
623 72
5 2 40 0 0 4224 0 27 18 0 0 3
419 256
617 256
617 72
5 3 41 0 0 4224 0 26 18 0 0 3
419 179
611 179
611 72
5 4 42 0 0 4224 0 25 18 0 0 3
419 102
605 102
605 72
1 3 43 0 0 4224 0 3 28 0 0 4
47 349
324 349
324 353
352 353
4 3 44 0 0 8320 0 25 32 0 0 6
419 120
432 120
432 717
342 717
342 693
350 693
4 3 45 0 0 12416 0 32 31 0 0 5
416 693
421 693
421 635
350 635
350 606
4 3 46 0 0 12416 0 31 30 0 0 6
416 606
421 606
421 530
338 530
338 516
351 516
4 3 47 0 0 12416 0 30 29 0 0 5
417 516
423 516
423 458
351 458
351 433
4 3 48 0 0 12416 0 26 25 0 0 6
419 197
423 197
423 140
345 140
345 120
353 120
4 3 49 0 0 12416 0 27 26 0 0 6
419 274
423 274
423 218
345 218
345 197
353 197
4 3 50 0 0 12416 0 28 27 0 0 6
418 353
423 353
423 288
345 288
345 274
353 274
4 8 18 0 0 0 0 21 21 0 0 6
93 595
89 595
89 610
171 610
171 595
163 595
4 8 22 0 0 0 0 22 22 0 0 6
95 496
91 496
91 511
173 511
173 496
165 496
1 2 51 0 0 8192 0 4 21 0 0 4
46 540
80 540
80 577
99 577
1 1 51 0 0 4224 0 4 21 0 0 4
46 540
85 540
85 568
99 568
1 2 52 0 0 8192 0 6 22 0 0 4
46 441
82 441
82 478
101 478
1 1 52 0 0 4224 0 6 22 0 0 4
46 441
87 441
87 469
101 469
1 3 53 0 0 4224 0 5 21 0 0 4
47 585
85 585
85 586
93 586
1 3 54 0 0 4224 0 7 22 0 0 4
44 489
87 489
87 487
95 487
1 1 55 0 0 4224 0 24 32 0 0 3
211 77
211 675
350 675
2 1 56 0 0 4224 0 24 31 0 0 3
205 77
205 588
350 588
3 1 57 0 0 4224 0 24 30 0 0 3
199 77
199 498
351 498
4 1 58 0 0 4224 0 24 29 0 0 3
193 77
193 415
351 415
1 1 59 0 0 4224 0 23 28 0 0 3
261 76
261 335
352 335
2 1 60 0 0 4224 0 23 27 0 0 3
255 76
255 256
353 256
3 1 61 0 0 8320 0 23 26 0 0 3
249 76
249 179
353 179
4 1 62 0 0 8320 0 23 25 0 0 3
243 76
243 102
353 102
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
