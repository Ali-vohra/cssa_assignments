CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 80 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
30
13 Logic Switch~
5 408 243 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89861e-315 0
0
13 Logic Switch~
5 28 387 0 1 11
0 25
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89861e-315 0
0
13 Logic Switch~
5 28 437 0 1 11
0 26
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89861e-315 0
0
13 Logic Switch~
5 159 574 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
43355.3 0
0
13 Logic Switch~
5 116 575 0 10 11
0 35 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8157 0 0
2
43355.3 1
0
13 Logic Switch~
5 28 488 0 1 11
0 27
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
5.89861e-315 5.26354e-315
0
9 Inverter~
13 397 381 0 2 22
0 5 4
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U10F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
8901 0 0
2
5.89861e-315 0
0
9 2-In AND~
219 405 428 0 3 22
0 4 3 2
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U15C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
7361 0 0
2
5.89861e-315 0
0
8 2-In OR~
219 395 316 0 3 22
0 7 6 3
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U16A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
4747 0 0
2
5.89861e-315 0
0
9 2-In AND~
219 404 141 0 3 22
0 9 8 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U15B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
972 0 0
2
5.89861e-315 0
0
9 2-In AND~
219 404 86 0 3 22
0 9 10 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U15A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3472 0 0
2
5.89861e-315 0
0
12 Hex Display~
7 665 40 0 18 19
10 12 13 14 15 0 0 0 0 0
0 1 1 1 1 0 1 1 9
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
9998 0 0
2
5.89861e-315 0
0
6 74LS90
107 124 470 0 10 21
0 25 25 26 26 27 21 24 23 22
21
0
0 0 4848 0
6 74LS90
-21 -51 21 -43
2 U5
-7 -52 7 -44
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
3536 0 0
2
5.89861e-315 0
0
9 Inverter~
13 248 470 0 2 22
0 24 39
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U10E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
4597 0 0
2
43355.3 2
0
9 Inverter~
13 247 686 0 2 22
0 21 36
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U10D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
3835 0 0
2
43355.3 3
0
9 Inverter~
13 246 611 0 2 22
0 22 37
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U10C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3670 0 0
2
43355.3 4
0
9 Inverter~
13 248 537 0 2 22
0 23 38
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U10B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
5616 0 0
2
43355.3 5
0
8 Hex Key~
166 118 46 0 11 12
0 43 44 45 46 0 0 0 0 0
0 48
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
9323 0 0
2
5.89861e-315 5.3568e-315
0
2 FA
94 302 111 0 5 11
0 46 31 40 5 9
2 FA
1 0 688 0
0
2 U1
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 1 0 0 0
1 U
317 0 0
2
5.89861e-315 5.36716e-315
0
2 FA
94 302 195 0 5 11
0 45 30 41 40 10
2 FA
2 0 688 0
0
2 U2
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 1 0 0 0
1 U
3108 0 0
2
5.89861e-315 5.37752e-315
0
2 FA
94 302 282 0 5 11
0 44 29 42 41 8
2 FA
3 0 688 0
0
2 U3
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 1 0 0 0
1 U
4299 0 0
2
5.89861e-315 5.38788e-315
0
2 FA
94 302 369 0 5 11
0 43 28 25 42 20
2 FA
4 0 688 0
0
2 U4
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 1 0 0 0
1 U
9672 0 0
2
5.89861e-315 5.39306e-315
0
2 FA
94 302 470 0 5 11
0 39 11 32 59 31
2 FA
5 0 688 0
0
2 U6
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 1 0 0 0
1 U
7876 0 0
2
43355.3 6
0
2 FA
94 301 537 0 5 11
0 38 11 33 32 30
2 FA
6 0 688 0
0
2 U7
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 1 0 0 0
1 U
6369 0 0
2
43355.3 7
0
2 FA
94 299 611 0 5 11
0 37 11 34 33 29
2 FA
7 0 688 0
0
2 U8
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 1 0 0 0
1 U
9172 0 0
2
43355.3 8
0
2 FA
94 298 686 0 5 11
0 36 35 11 34 28
2 FA
8 0 688 0
0
2 U9
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 1 0 0 0
1 U
7100 0 0
2
43355.3 9
0
2 FA
94 496 111 0 5 11
0 9 2 16 72 15
2 FA
9 0 688 0
0
3 U11
-11 -29 10 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 1 0 0 0
1 U
3820 0 0
2
5.89859e-315 0
0
2 FA
94 496 195 0 5 11
0 10 19 17 16 14
2 FA
10 0 688 0
0
3 U12
-11 -29 10 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 1 0 0 0
1 U
7678 0 0
2
5.89859e-315 0
0
2 FA
94 495 282 0 5 11
0 8 2 18 17 13
2 FA
11 0 688 0
0
3 U13
-11 -29 10 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 1 0 0 0
1 U
961 0 0
2
5.89859e-315 0
0
2 FA
94 496 369 0 5 11
0 20 19 19 18 12
2 FA
12 0 688 0
0
3 U14
-11 -29 10 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 1 0 0 0
1 U
3178 0 0
2
5.89859e-315 0
0
59
3 2 2 0 0 8192 0 8 29 0 0 4
426 428
449 428
449 291
462 291
3 2 2 0 0 8320 0 8 27 0 0 4
426 428
435 428
435 120
463 120
3 2 3 0 0 8320 0 9 8 0 0 6
428 316
452 316
452 448
373 448
373 437
381 437
2 1 4 0 0 12416 0 7 8 0 0 6
418 381
430 381
430 408
373 408
373 419
381 419
4 1 5 0 0 8320 0 19 7 0 0 4
335 129
364 129
364 381
382 381
3 2 6 0 0 8320 0 11 9 0 0 6
425 86
437 86
437 336
374 336
374 325
382 325
3 1 7 0 0 8320 0 10 9 0 0 6
425 141
432 141
432 296
374 296
374 307
382 307
5 2 8 0 0 8320 0 21 10 0 0 4
335 282
371 282
371 150
380 150
5 1 9 0 0 4096 0 19 10 0 0 4
335 111
361 111
361 132
380 132
5 2 10 0 0 8192 0 20 11 0 0 4
335 195
367 195
367 95
380 95
5 1 9 0 0 4096 0 19 11 0 0 4
335 111
372 111
372 77
380 77
0 3 11 0 0 8192 0 0 26 38 0 4
171 619
227 619
227 704
265 704
5 1 12 0 0 8320 0 30 12 0 0 3
529 369
674 369
674 64
5 2 13 0 0 8320 0 29 12 0 0 3
528 282
668 282
668 64
5 3 14 0 0 4224 0 28 12 0 0 3
529 195
662 195
662 64
5 4 15 0 0 4224 0 27 12 0 0 3
529 111
656 111
656 64
4 3 16 0 0 12416 0 28 27 0 0 5
529 213
533 213
533 153
463 153
463 129
4 3 17 0 0 12416 0 29 28 0 0 6
528 300
533 300
533 227
445 227
445 213
463 213
4 3 18 0 0 12416 0 30 29 0 0 6
529 387
532 387
532 314
454 314
454 300
462 300
1 3 19 0 0 8320 0 1 30 0 0 4
420 243
440 243
440 387
463 387
1 2 19 0 0 0 0 1 30 0 0 4
420 243
445 243
445 378
463 378
1 2 19 0 0 0 0 1 28 0 0 4
420 243
455 243
455 204
463 204
5 1 20 0 0 4224 0 22 30 0 0 2
335 369
463 369
5 1 8 0 0 0 0 21 29 0 0 2
335 282
462 282
5 1 10 0 0 4224 0 20 28 0 0 2
335 195
463 195
5 1 9 0 0 4224 0 19 27 0 0 2
335 111
463 111
10 1 21 0 0 8320 0 13 15 0 0 4
156 497
214 497
214 686
232 686
9 1 22 0 0 8320 0 13 16 0 0 4
156 479
223 479
223 611
231 611
8 1 23 0 0 8320 0 13 17 0 0 4
156 461
220 461
220 537
233 537
7 1 24 0 0 4224 0 13 14 0 0 4
156 443
225 443
225 470
233 470
1 3 25 0 0 4224 0 2 22 0 0 2
40 387
269 387
1 2 25 0 0 0 0 2 13 0 0 4
40 387
63 387
63 452
92 452
1 1 25 0 0 0 0 2 13 0 0 4
40 387
68 387
68 443
92 443
1 4 26 0 0 4096 0 3 13 0 0 4
40 437
73 437
73 470
92 470
1 3 26 0 0 4224 0 3 13 0 0 4
40 437
78 437
78 461
92 461
10 6 21 0 0 0 0 13 13 0 0 6
156 497
160 497
160 512
78 512
78 497
86 497
1 5 27 0 0 4224 0 6 13 0 0 2
40 488
86 488
1 2 11 0 0 8192 0 4 25 0 0 3
171 574
171 620
266 620
1 2 11 0 0 8192 0 4 24 0 0 3
171 574
171 546
268 546
1 2 11 0 0 8320 0 4 23 0 0 3
171 574
171 479
269 479
5 2 28 0 0 8320 0 26 22 0 0 6
331 686
359 686
359 345
261 345
261 378
269 378
5 2 29 0 0 8320 0 25 21 0 0 6
332 611
349 611
349 258
261 258
261 291
269 291
5 2 30 0 0 8320 0 24 20 0 0 6
334 537
344 537
344 227
261 227
261 204
269 204
5 2 31 0 0 8320 0 23 19 0 0 6
335 470
339 470
339 87
261 87
261 120
269 120
4 3 32 0 0 12416 0 24 23 0 0 6
334 555
339 555
339 502
261 502
261 488
269 488
4 3 33 0 0 12416 0 25 24 0 0 6
332 629
338 629
338 569
260 569
260 555
268 555
4 3 34 0 0 12416 0 26 25 0 0 6
331 704
336 704
336 643
258 643
258 629
266 629
1 2 35 0 0 8320 0 5 26 0 0 3
128 575
128 695
265 695
1 2 36 0 0 4224 0 26 15 0 0 2
265 686
268 686
1 2 37 0 0 4224 0 25 16 0 0 2
266 611
267 611
1 2 38 0 0 4224 0 24 17 0 0 2
268 537
269 537
2 1 39 0 0 4224 0 14 23 0 0 4
269 470
271 470
271 470
269 470
4 3 40 0 0 12416 0 20 19 0 0 5
335 213
353 213
353 156
269 156
269 129
4 3 41 0 0 12416 0 21 20 0 0 5
335 300
353 300
353 242
269 242
269 213
4 3 42 0 0 12416 0 22 21 0 0 5
335 387
353 387
353 329
269 329
269 300
1 1 43 0 0 4224 0 18 22 0 0 3
127 70
127 369
269 369
2 1 44 0 0 4224 0 18 21 0 0 3
121 70
121 282
269 282
3 1 45 0 0 8320 0 18 20 0 0 3
115 70
115 195
269 195
4 1 46 0 0 8320 0 18 19 0 0 3
109 70
109 111
269 111
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
