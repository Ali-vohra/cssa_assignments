CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
100 20 5 120 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
15
13 Logic Switch~
5 680 271 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43329.9 0
0
13 Logic Switch~
5 115 277 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
43329.9 0
0
12 Hex Display~
7 876 64 0 16 19
10 10 11 12 13 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3124 0 0
2
43329.9 0
0
12 Hex Display~
7 608 69 0 16 19
10 6 7 8 9 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3421 0 0
2
43329.9 0
0
12 Hex Display~
7 328 76 0 16 19
10 2 3 4 5 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
8157 0 0
2
43329.9 0
0
8 2-In OR~
219 421 158 0 3 22
0 17 18 16
0
0 0 624 180
6 74LS32
-21 -24 21 -16
3 U6A
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
5572 0 0
2
43329.9 0
0
5 4073~
219 230 162 0 4 22
0 21 20 19 18
0
0 0 624 180
4 4073
-7 -24 21 -16
3 U5A
-13 -25 8 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 2 0
1 U
8901 0 0
2
43329.9 0
0
9 2-In AND~
219 229 218 0 3 22
0 3 3 21
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U4D
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
7361 0 0
2
43329.9 0
0
9 2-In AND~
219 489 196 0 3 22
0 7 6 20
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U4C
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
4747 0 0
2
43329.9 0
0
9 2-In AND~
219 776 219 0 3 22
0 13 10 19
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U4B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
972 0 0
2
43329.9 0
0
9 2-In AND~
219 491 248 0 3 22
0 6 9 17
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U4A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3472 0 0
2
43329.9 0
0
7 Pulser~
4 643 444 0 10 12
0 23 24 22 25 0 0 5 5 3
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
9998 0 0
2
43329.9 0
0
6 74LS90
107 774 297 0 10 21
0 14 14 18 18 22 10 13 12 11
10
0
0 0 4848 0
6 74LS90
-21 -51 21 -43
2 U3
-7 -52 7 -44
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 0 0 0 0
1 U
3536 0 0
2
43329.9 0
0
6 74LS93
109 490 309 0 8 17
0 16 16 13 6 9 8 7 6
0
0 0 4848 0
6 74LS93
-21 -35 21 -27
2 U2
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 0 0 0 0
1 U
4597 0 0
2
43329.9 0
0
6 74LS90
107 227 301 0 10 21
0 15 15 18 18 9 2 5 4 3
2
0
0 0 4848 0
6 74LS90
-21 -51 21 -43
2 U1
-7 -52 7 -44
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 0 0 0 0
1 U
3835 0 0
2
43329.9 0
0
41
10 1 2 0 0 8320 0 15 5 0 0 3
259 328
337 328
337 100
9 2 3 0 0 8320 0 15 5 0 0 3
259 310
331 310
331 100
8 3 4 0 0 8320 0 15 5 0 0 3
259 292
325 292
325 100
7 4 5 0 0 8320 0 15 5 0 0 3
259 274
319 274
319 100
8 1 6 0 0 8320 0 14 4 0 0 3
522 327
617 327
617 93
7 2 7 0 0 8320 0 14 4 0 0 3
522 318
611 318
611 93
6 3 8 0 0 8320 0 14 4 0 0 3
522 309
605 309
605 93
5 4 9 0 0 8192 0 14 4 0 0 3
522 300
599 300
599 93
10 1 10 0 0 8320 0 13 3 0 0 3
806 324
885 324
885 88
9 2 11 0 0 8320 0 13 3 0 0 3
806 306
879 306
879 88
8 3 12 0 0 8320 0 13 3 0 0 3
806 288
873 288
873 88
7 4 13 0 0 8192 0 13 3 0 0 3
806 270
867 270
867 88
1 2 14 0 0 4096 0 1 13 0 0 4
692 271
723 271
723 279
742 279
1 1 14 0 0 4224 0 1 13 0 0 4
692 271
728 271
728 270
742 270
1 2 15 0 0 4096 0 2 15 0 0 4
127 277
161 277
161 283
195 283
1 1 15 0 0 4224 0 2 15 0 0 4
127 277
166 277
166 274
195 274
3 2 16 0 0 4224 0 6 14 0 0 3
394 158
394 309
458 309
3 1 16 0 0 0 0 6 14 0 0 4
394 158
382 158
382 300
458 300
3 1 17 0 0 8320 0 11 6 0 0 4
464 248
450 248
450 167
440 167
4 2 18 0 0 12288 0 7 6 0 0 8
203 162
194 162
194 245
387 245
387 274
445 274
445 149
440 149
4 4 18 0 0 12416 0 7 13 0 0 6
203 162
170 162
170 363
718 363
718 297
742 297
4 3 18 0 0 0 0 7 13 0 0 6
203 162
185 162
185 358
723 358
723 288
742 288
4 4 18 0 0 0 0 7 15 0 0 4
203 162
176 162
176 301
195 301
4 3 18 0 0 0 0 7 15 0 0 4
203 162
181 162
181 292
195 292
3 3 19 0 0 4224 0 10 7 0 0 4
749 219
268 219
268 153
248 153
3 2 20 0 0 4224 0 9 7 0 0 4
462 196
263 196
263 162
248 162
3 1 21 0 0 8320 0 8 7 0 0 6
202 218
201 218
201 142
258 142
258 171
248 171
2 9 3 0 0 0 0 8 15 0 0 4
247 209
272 209
272 310
259 310
1 9 3 0 0 0 0 8 15 0 0 4
247 227
267 227
267 310
259 310
2 8 6 0 0 0 0 9 14 0 0 4
507 187
545 187
545 327
522 327
1 7 7 0 0 0 0 9 14 0 0 4
507 205
540 205
540 318
522 318
2 10 10 0 0 0 0 10 13 0 0 4
794 210
819 210
819 324
806 324
1 7 13 0 0 0 0 10 13 0 0 4
794 228
814 228
814 270
806 270
1 8 6 0 0 0 0 11 14 0 0 4
509 257
535 257
535 327
522 327
2 5 9 0 0 0 0 11 14 0 0 4
509 239
530 239
530 300
522 300
10 6 2 0 0 0 0 15 15 0 0 6
259 328
263 328
263 343
176 343
176 328
189 328
5 5 9 0 0 12416 0 14 15 0 0 6
522 300
526 300
526 352
181 352
181 319
189 319
4 8 6 0 0 0 0 14 14 0 0 6
452 327
448 327
448 347
530 347
530 327
522 327
7 3 13 0 0 12416 0 13 14 0 0 6
806 270
810 270
810 342
444 342
444 318
452 318
6 10 10 0 0 0 0 13 13 0 0 6
736 324
732 324
732 339
814 339
814 324
806 324
3 5 22 0 0 8320 0 12 13 0 0 4
667 435
728 435
728 315
736 315
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
430 494 605 518
437 500 597 516
20 3 BIT COUNTER(COMB.)
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
