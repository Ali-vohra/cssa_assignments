CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 568 528 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V5
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43382.9 0
0
13 Logic Switch~
5 517 530 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V4
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
391 0 0
2
43382.9 0
0
13 Logic Switch~
5 471 530 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V3
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3124 0 0
2
43382.9 0
0
13 Logic Switch~
5 190 204 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3421 0 0
2
43382.9 0
0
13 Logic Switch~
5 191 164 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8157 0 0
2
43382.9 0
0
14 Logic Display~
6 755 263 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5572 0 0
2
43382.9 0
0
9 Inverter~
13 337 392 0 2 22
0 7 6
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
8901 0 0
2
43382.9 0
0
9 2-In AND~
219 346 319 0 3 22
0 7 9 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
7361 0 0
2
43382.9 0
0
9 2-In XOR~
219 342 248 0 3 22
0 7 9 10
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U3A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
4747 0 0
2
43382.9 0
0
8 2-In OR~
219 341 173 0 3 22
0 7 9 11
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
972 0 0
2
43382.9 0
0
8 4x1 MUX~
94 470 285 0 8 17
0 11 10 8 6 5 3 4 2
7 4x1 MUX
1 0 560 0
0
2 U1
1 -68 15 -60
0
0
0
0
0
0
17

0 3 4 5 6 9 12 13 16 3
4 5 6 9 12 13 16 0
0 0 0 0 0 0 0 0
1 U
3472 0 0
2
43361.9 0
0
15
1 8 2 0 0 4224 0 1 11 0 0 3
569 515
569 250
519 250
1 6 3 0 0 4224 0 2 11 0 0 5
518 517
518 353
532 353
532 296
519 296
1 7 4 0 0 4224 0 3 11 0 0 5
472 517
472 348
527 348
527 285
519 285
5 1 5 0 0 4224 0 11 6 0 0 3
519 331
755 331
755 281
2 4 6 0 0 8320 0 7 11 0 0 4
358 392
424 392
424 308
437 308
0 1 7 0 0 4224 0 0 7 9 0 3
261 164
261 392
322 392
3 3 8 0 0 4224 0 8 11 0 0 4
367 319
429 319
429 296
437 296
1 2 9 0 0 8320 0 4 8 0 0 4
202 204
271 204
271 328
322 328
1 1 7 0 0 0 0 5 8 0 0 4
203 164
276 164
276 310
322 310
3 2 10 0 0 4224 0 9 11 0 0 4
375 248
424 248
424 285
437 285
1 2 9 0 0 0 0 4 9 0 0 4
202 204
282 204
282 257
326 257
1 1 7 0 0 0 0 5 9 0 0 4
203 164
287 164
287 239
326 239
3 1 11 0 0 8320 0 10 11 0 0 4
374 173
429 173
429 274
437 274
1 2 9 0 0 0 0 4 10 0 0 4
202 204
292 204
292 182
328 182
1 1 7 0 0 0 0 5 10 0 0 2
203 164
328 164
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
776 251 805 275
786 259 794 275
1 F
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
557 564 586 588
567 572 575 588
1 E
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
503 564 540 588
513 572 529 588
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
456 564 493 588
466 572 482 588
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
133 184 170 208
143 192 159 208
2 B0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
133 143 170 167
143 151 159 167
2 A0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
