CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
160 250 7 140 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
14
13 Logic Switch~
5 646 311 0 1 11
0 14
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 388 317 0 1 11
0 15
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 177 318 0 1 11
0 16
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89855e-315 0
0
12 Hex Display~
7 738 70 0 16 19
10 2 3 4 5 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3421 0 0
2
5.89855e-315 0
0
12 Hex Display~
7 508 78 0 18 19
10 6 7 8 9 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
8157 0 0
2
5.89855e-315 0
0
12 Hex Display~
7 279 84 0 16 19
10 10 11 12 13 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
5572 0 0
2
5.89855e-315 0
0
5 4073~
219 509 173 0 4 22
0 20 19 18 17
0
0 0 608 180
4 4073
-7 -24 21 -16
3 U5A
-13 -25 8 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 2 0
1 U
8901 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 283 248 0 3 22
0 11 11 20
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U4C
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
7361 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 512 247 0 3 22
0 7 6 19
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U4B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
4747 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 744 245 0 3 22
0 5 2 18
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U4A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
972 0 0
2
5.89855e-315 0
0
7 Pulser~
4 665 429 0 10 12
0 22 23 21 24 0 0 5 5 2
7
0
0 0 4640 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3472 0 0
2
5.89855e-315 0
0
6 74LS90
107 744 338 0 10 21
0 14 14 17 17 21 2 5 4 3
2
0
0 0 4832 0
6 74LS90
-21 -51 21 -43
2 U3
-7 -52 7 -44
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
9998 0 0
2
5.89855e-315 0
0
6 74LS90
107 508 338 0 10 21
0 15 15 17 17 5 6 9 8 7
6
0
0 0 4832 0
6 74LS90
-21 -51 21 -43
2 U2
-7 -52 7 -44
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
3536 0 0
2
5.89855e-315 0
0
6 74LS90
107 280 339 0 10 21
0 16 16 17 17 9 10 13 12 11
10
0
0 0 4832 0
6 74LS90
-21 -51 21 -43
2 U1
-7 -52 7 -44
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
4597 0 0
2
5.89855e-315 0
0
39
10 1 2 0 0 8320 0 12 4 0 0 5
776 365
810 365
810 117
747 117
747 94
9 2 3 0 0 8320 0 12 4 0 0 5
776 347
805 347
805 112
741 112
741 94
8 3 4 0 0 8320 0 12 4 0 0 5
776 329
800 329
800 107
735 107
735 94
7 4 5 0 0 8192 0 12 4 0 0 5
776 311
795 311
795 102
729 102
729 94
10 1 6 0 0 8320 0 13 5 0 0 5
540 365
574 365
574 125
517 125
517 102
9 2 7 0 0 8320 0 13 5 0 0 5
540 347
569 347
569 120
511 120
511 102
8 3 8 0 0 8320 0 13 5 0 0 5
540 329
564 329
564 115
505 115
505 102
7 4 9 0 0 8192 0 13 5 0 0 5
540 311
559 311
559 110
499 110
499 102
10 1 10 0 0 8320 0 14 6 0 0 5
312 366
341 366
341 131
288 131
288 108
9 2 11 0 0 8320 0 14 6 0 0 5
312 348
336 348
336 126
282 126
282 108
8 3 12 0 0 8320 0 14 6 0 0 5
312 330
331 330
331 121
276 121
276 108
7 4 13 0 0 8320 0 14 6 0 0 5
312 312
326 312
326 116
270 116
270 108
1 2 14 0 0 4096 0 1 12 0 0 4
658 311
698 311
698 320
712 320
1 1 14 0 0 4224 0 1 12 0 0 2
658 311
712 311
1 2 15 0 0 4096 0 2 13 0 0 4
400 317
442 317
442 320
476 320
1 1 15 0 0 4224 0 2 13 0 0 4
400 317
447 317
447 311
476 311
1 2 16 0 0 4096 0 3 14 0 0 4
189 318
219 318
219 321
248 321
1 1 16 0 0 4224 0 3 14 0 0 4
189 318
224 318
224 312
248 312
4 4 17 0 0 12288 0 7 12 0 0 6
482 173
451 173
451 400
683 400
683 338
712 338
4 3 17 0 0 0 0 7 12 0 0 6
482 173
466 173
466 395
688 395
688 329
712 329
4 4 17 0 0 0 0 7 13 0 0 4
482 173
457 173
457 338
476 338
4 3 17 0 0 0 0 7 13 0 0 4
482 173
462 173
462 329
476 329
4 4 17 0 0 4224 0 7 14 0 0 4
482 173
229 173
229 339
248 339
4 3 17 0 0 0 0 7 14 0 0 4
482 173
234 173
234 330
248 330
3 3 18 0 0 4224 0 10 7 0 0 4
717 245
547 245
547 164
527 164
3 2 19 0 0 8320 0 9 7 0 0 6
485 247
480 247
480 148
542 148
542 173
527 173
3 1 20 0 0 12416 0 8 7 0 0 6
256 248
254 248
254 153
537 153
537 182
527 182
9 2 11 0 0 0 0 14 8 0 0 4
312 348
321 348
321 239
301 239
9 1 11 0 0 0 0 14 8 0 0 4
312 348
316 348
316 257
301 257
10 2 6 0 0 0 0 13 9 0 0 4
540 365
554 365
554 238
530 238
9 1 7 0 0 0 0 13 9 0 0 4
540 347
544 347
544 256
530 256
10 2 2 0 0 0 0 12 10 0 0 4
776 365
790 365
790 236
762 236
7 1 5 0 0 0 0 12 10 0 0 4
776 311
780 311
780 254
762 254
10 6 10 0 0 0 0 14 14 0 0 6
312 366
316 366
316 381
229 381
229 366
242 366
7 5 9 0 0 12416 0 13 14 0 0 6
540 311
549 311
549 390
234 390
234 357
242 357
10 6 6 0 0 0 0 13 13 0 0 6
540 365
544 365
544 380
457 380
457 365
470 365
7 5 5 0 0 12416 0 12 13 0 0 6
776 311
785 311
785 385
462 385
462 356
470 356
10 6 2 0 0 0 0 12 12 0 0 6
776 365
780 365
780 380
693 380
693 365
706 365
3 5 21 0 0 8320 0 11 12 0 0 4
689 420
700 420
700 356
706 356
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
429 457 612 481
436 463 604 479
21 3 BIT COUNTER IC 7490
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
