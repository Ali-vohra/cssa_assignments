CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
25
13 Logic Switch~
5 788 357 0 1 11
0 7
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 543 360 0 1 11
0 19
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 161 230 0 1 11
0 20
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 163 424 0 10 11
0 39 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
5.89855e-315 0
0
12 Hex Display~
7 1108 138 0 16 19
10 2 3 4 5 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
8157 0 0
2
5.89855e-315 0
0
9 Inverter~
13 703 491 0 2 22
0 12 6
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
5572 0 0
2
5.89855e-315 0
0
5 4030~
219 878 495 0 3 22
0 13 6 8
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U8D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 4 0
1 U
8901 0 0
2
5.89855e-315 0
0
5 4030~
219 878 445 0 3 22
0 14 6 9
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U8C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 4 0
1 U
7361 0 0
2
5.89855e-315 0
0
5 4030~
219 878 396 0 3 22
0 15 6 10
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U8B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 4 0
1 U
4747 0 0
2
5.89855e-315 0
0
5 4030~
219 877 352 0 3 22
0 16 6 11
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U8A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
972 0 0
2
5.89855e-315 0
0
6 74LS83
105 966 268 0 14 29
0 6 7 6 7 11 10 9 8 6
5 4 3 2 44
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U7
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
3472 0 0
2
5.89855e-315 0
0
14 Logic Display~
6 669 163 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9998 0 0
2
5.89855e-315 0
0
14 Logic Display~
6 440 356 0 1 2
10 18
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3536 0 0
2
5.89855e-315 0
0
8 3-In OR~
219 657 421 0 4 22
0 21 17 22 12
0
0 0 608 270
4 4075
-14 -24 14 -16
3 U6A
28 -7 49 1
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 3 0
1 U
4597 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 694 361 0 3 22
0 23 24 21
0
0 0 608 270
6 74LS08
-21 -24 21 -16
3 U5B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3835 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 619 361 0 3 22
0 25 24 22
0
0 0 608 270
6 74LS08
-21 -24 21 -16
3 U5A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3670 0 0
2
5.89855e-315 0
0
6 74LS83
105 788 272 0 14 29
0 24 25 23 26 20 12 12 20 19
16 15 14 13 45
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U4
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
5616 0 0
2
5.89855e-315 0
0
8 Hex Key~
166 393 98 0 11 12
0 27 28 29 30 0 0 0 0 0
9 57
0
0 0 4640 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
9323 0 0
2
5.89855e-315 0
0
6 74LS83
105 544 275 0 14 29
0 30 29 28 27 34 33 32 31 20
24 25 23 26 17
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U3
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
317 0 0
2
5.89855e-315 0
0
8 Hex Key~
166 86 104 0 11 12
0 35 36 37 38 0 0 0 0 0
9 57
0
0 0 4640 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3108 0 0
2
5.89855e-315 0
0
9 Inverter~
13 161 376 0 2 22
0 35 40
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
4299 0 0
2
5.89855e-315 0
0
9 Inverter~
13 159 342 0 2 22
0 36 41
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
9672 0 0
2
5.89855e-315 0
0
9 Inverter~
13 158 307 0 2 22
0 37 42
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
7876 0 0
2
5.89855e-315 0
0
9 Inverter~
13 159 272 0 2 22
0 38 43
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
6369 0 0
2
5.89855e-315 0
0
6 74LS83
105 333 277 0 14 29
0 39 20 39 20 43 42 41 40 39
34 33 32 31 18
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
9172 0 0
2
5.89855e-315 0
0
62
13 1 2 0 0 8320 0 11 5 0 0 3
998 286
1117 286
1117 162
12 2 3 0 0 8320 0 11 5 0 0 3
998 277
1111 277
1111 162
11 3 4 0 0 4224 0 11 5 0 0 3
998 268
1105 268
1105 162
10 4 5 0 0 4224 0 11 5 0 0 3
998 259
1099 259
1099 162
2 9 6 0 0 8192 0 6 11 0 0 4
724 491
826 491
826 313
934 313
1 4 7 0 0 12288 0 1 11 0 0 4
800 357
827 357
827 259
934 259
1 2 7 0 0 8320 0 1 11 0 0 4
800 357
832 357
832 241
934 241
2 3 6 0 0 8192 0 6 11 0 0 4
724 491
836 491
836 250
934 250
2 1 6 0 0 8320 0 6 11 0 0 4
724 491
856 491
856 232
934 232
3 8 8 0 0 8320 0 7 11 0 0 4
911 495
916 495
916 295
934 295
3 7 9 0 0 8320 0 8 11 0 0 4
911 445
916 445
916 286
934 286
3 6 10 0 0 8320 0 9 11 0 0 4
911 396
921 396
921 277
934 277
3 5 11 0 0 8320 0 10 11 0 0 4
910 352
926 352
926 268
934 268
2 2 6 0 0 0 0 6 7 0 0 4
724 491
839 491
839 504
862 504
2 2 6 0 0 0 0 6 8 0 0 4
724 491
844 491
844 454
862 454
2 2 6 0 0 0 0 6 9 0 0 4
724 491
849 491
849 405
862 405
2 2 6 0 0 0 0 6 10 0 0 4
724 491
853 491
853 361
861 361
4 1 12 0 0 4096 0 14 6 0 0 3
660 451
660 491
688 491
13 1 13 0 0 8320 0 17 7 0 0 4
820 290
839 290
839 486
862 486
12 1 14 0 0 8320 0 17 8 0 0 4
820 281
844 281
844 436
862 436
11 1 15 0 0 8320 0 17 9 0 0 4
820 272
849 272
849 387
862 387
10 1 16 0 0 8320 0 17 10 0 0 4
820 263
853 263
853 343
861 343
14 1 17 0 0 8320 0 19 12 0 0 3
576 320
669 320
669 181
14 1 18 0 0 4224 0 25 13 0 0 5
365 322
427 322
427 382
440 382
440 374
1 9 19 0 0 12416 0 2 17 0 0 4
555 360
598 360
598 317
756 317
1 8 20 0 0 12416 0 3 17 0 0 6
173 230
267 230
267 394
738 394
738 299
756 299
1 5 20 0 0 0 0 3 17 0 0 6
173 230
282 230
282 219
728 219
728 272
756 272
4 7 12 0 0 12288 0 14 17 0 0 5
660 451
660 453
743 453
743 290
756 290
4 6 12 0 0 12416 0 14 17 0 0 5
660 451
660 448
748 448
748 281
756 281
14 2 17 0 0 0 0 19 14 0 0 3
576 320
660 320
660 406
3 1 21 0 0 8320 0 15 14 0 0 4
692 384
692 390
669 390
669 405
3 3 22 0 0 8320 0 16 14 0 0 4
617 384
617 390
651 390
651 405
12 1 23 0 0 4096 0 19 15 0 0 3
576 284
701 284
701 339
10 2 24 0 0 4096 0 19 15 0 0 3
576 266
683 266
683 339
11 1 25 0 0 8192 0 19 16 0 0 3
576 275
626 275
626 339
10 2 24 0 0 0 0 19 16 0 0 3
576 266
608 266
608 339
13 4 26 0 0 4224 0 19 17 0 0 4
576 293
733 293
733 263
756 263
12 3 23 0 0 4224 0 19 17 0 0 4
576 284
738 284
738 254
756 254
11 2 25 0 0 4224 0 19 17 0 0 4
576 275
743 275
743 245
756 245
10 1 24 0 0 4224 0 19 17 0 0 4
576 266
748 266
748 236
756 236
1 9 20 0 0 0 0 3 19 0 0 6
173 230
297 230
297 337
504 337
504 320
512 320
1 4 27 0 0 4224 0 18 19 0 0 3
402 122
402 266
512 266
2 3 28 0 0 4224 0 18 19 0 0 3
396 122
396 257
512 257
3 2 29 0 0 4224 0 18 19 0 0 3
390 122
390 248
512 248
4 1 30 0 0 8320 0 18 19 0 0 3
384 122
384 239
512 239
13 8 31 0 0 4224 0 25 19 0 0 4
365 295
504 295
504 302
512 302
12 7 32 0 0 4224 0 25 19 0 0 4
365 286
504 286
504 293
512 293
11 6 33 0 0 4224 0 25 19 0 0 4
365 277
504 277
504 284
512 284
10 5 34 0 0 4224 0 25 19 0 0 4
365 268
504 268
504 275
512 275
1 1 35 0 0 4224 0 20 21 0 0 3
95 128
95 376
146 376
2 1 36 0 0 4224 0 20 22 0 0 3
89 128
89 342
144 342
3 1 37 0 0 4224 0 20 23 0 0 3
83 128
83 307
143 307
4 1 38 0 0 4224 0 20 24 0 0 3
77 128
77 272
144 272
1 4 20 0 0 0 0 3 25 0 0 4
173 230
288 230
288 268
301 268
1 2 20 0 0 0 0 3 25 0 0 4
173 230
293 230
293 250
301 250
1 3 39 0 0 8192 0 4 25 0 0 4
175 424
273 424
273 259
301 259
1 1 39 0 0 8320 0 4 25 0 0 4
175 424
278 424
278 241
301 241
1 9 39 0 0 0 0 4 25 0 0 4
175 424
293 424
293 322
301 322
2 8 40 0 0 4224 0 21 25 0 0 4
182 376
283 376
283 304
301 304
2 7 41 0 0 4224 0 22 25 0 0 4
180 342
288 342
288 295
301 295
2 6 42 0 0 4224 0 23 25 0 0 4
179 307
293 307
293 286
301 286
2 5 43 0 0 4224 0 24 25 0 0 4
180 272
293 272
293 277
301 277
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
455 541 644 565
465 549 633 565
21 BCD SUBTRACTOR (10'S)
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
