CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
16
13 Logic Switch~
5 71 94 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 69 228 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 70 177 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 72 51 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 352 398 0 3 22
0 4 3 2
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-13 -3 8 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
8157 0 0
2
43337.5 0
0
9 2-In XOR~
219 346 353 0 3 22
0 4 3 12
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U2B
-1 -3 20 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
5572 0 0
2
43337.5 0
0
9 2-In AND~
219 217 397 0 3 22
0 5 6 4
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-13 -3 8 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
8901 0 0
2
43337.5 0
0
9 2-In XOR~
219 212 351 0 3 22
0 6 5 7
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U2A
0 -2 21 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
7361 0 0
2
43337.5 0
0
14 Logic Display~
6 504 443 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4747 0 0
2
5.89859e-315 0
0
14 Logic Display~
6 416 445 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
972 0 0
2
5.89859e-315 0
0
14 Logic Display~
6 301 447 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3472 0 0
2
5.89859e-315 0
0
14 Logic Display~
6 159 450 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9998 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 350 278 0 3 22
0 8 9 3
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1D
-13 -12 8 -4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
3536 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 242 277 0 3 22
0 8 10 5
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1C
-12 -11 9 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
4597 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 202 277 0 3 22
0 11 9 6
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1B
-12 -11 9 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3835 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 133 276 0 3 22
0 11 10 13
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1A
-12 -11 9 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3670 0 0
2
5.89859e-315 0
0
24
3 1 2 0 0 4224 0 5 9 0 0 5
373 398
474 398
474 478
504 478
504 461
0 2 3 0 0 4096 0 0 5 5 0 3
301 362
301 407
328 407
1 0 4 0 0 4096 0 5 0 0 4 2
328 389
310 389
3 1 4 0 0 4224 0 7 6 0 0 4
238 397
310 397
310 344
330 344
3 2 3 0 0 12416 0 13 6 0 0 5
348 301
348 314
301 314
301 362
330 362
0 1 5 0 0 4096 0 0 7 10 0 3
185 360
185 388
193 388
0 2 6 0 0 4224 0 0 7 9 0 3
177 342
177 406
193 406
3 1 7 0 0 8320 0 8 11 0 0 5
245 351
275 351
275 479
301 479
301 465
3 1 6 0 0 0 0 15 8 0 0 5
200 300
200 313
177 313
177 342
196 342
3 2 5 0 0 8320 0 14 8 0 0 5
240 300
240 320
185 320
185 360
196 360
1 0 8 0 0 4096 0 13 0 0 20 2
357 256
357 177
2 0 9 0 0 4096 0 13 0 0 22 2
339 256
339 51
1 0 8 0 0 0 0 14 0 0 20 2
249 255
249 177
2 0 10 0 0 4096 0 14 0 0 21 2
231 255
231 94
1 0 11 0 0 4096 0 15 0 0 19 2
209 255
209 228
2 0 9 0 0 0 0 15 0 0 22 2
191 255
191 51
1 0 11 0 0 0 0 16 0 0 19 2
140 254
140 228
2 0 10 0 0 0 0 16 0 0 21 2
122 254
122 94
1 0 11 0 0 4224 0 2 0 0 0 2
81 228
523 228
1 0 8 0 0 4224 0 3 0 0 0 2
82 177
523 177
1 0 10 0 0 4224 0 1 0 0 0 2
83 94
524 94
1 0 9 0 0 4224 0 4 0 0 0 2
84 51
524 51
3 1 12 0 0 8320 0 6 10 0 0 5
379 353
394 353
394 478
416 478
416 463
3 1 13 0 0 4224 0 16 12 0 0 4
131 299
131 477
159 477
159 468
8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
18 32 55 56
28 40 44 56
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
16 75 53 99
26 83 42 99
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
15 156 52 180
25 164 41 180
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
14 204 51 228
24 212 40 228
2 B0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
141 501 178 525
151 509 167 525
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
284 500 321 524
294 508 310 524
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
398 501 435 525
408 509 424 525
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
490 501 527 525
500 509 516 525
2 S3
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
