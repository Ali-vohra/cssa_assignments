CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
20
13 Logic Switch~
5 585 233 0 1 11
0 6
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 344 287 0 1 11
0 17
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 143 427 0 1 11
0 30
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 139 228 0 10 11
0 31 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
5.89855e-315 0
0
12 Hex Display~
7 789 127 0 18 19
10 2 3 4 5 0 0 0 0 0
0 1 1 1 1 0 1 1 9
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
8157 0 0
2
5.89855e-315 0
0
9 Inverter~
13 512 370 0 2 22
0 7 12
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
5572 0 0
2
5.89855e-315 0
0
5 4030~
219 583 527 0 3 22
0 13 12 8
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U6D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 2 0
1 U
8901 0 0
2
5.89855e-315 0
0
5 4030~
219 582 474 0 3 22
0 14 12 9
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U6C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
7361 0 0
2
5.89855e-315 0
0
5 4030~
219 580 421 0 3 22
0 15 12 10
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U6B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
4747 0 0
2
5.89855e-315 0
0
5 4030~
219 579 367 0 3 22
0 16 12 11
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U6A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
972 0 0
2
5.89855e-315 0
0
6 74LS83
105 677 268 0 14 29
0 6 6 6 6 11 10 9 8 7
5 4 3 2 40
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U5
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
3472 0 0
2
5.89855e-315 0
0
6 74LS83
105 474 274 0 14 29
0 25 24 23 22 21 20 19 18 17
16 15 14 13 7
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U3
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
9998 0 0
2
5.89855e-315 0
0
9 Inverter~
13 330 584 0 2 22
0 26 18
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
3536 0 0
2
5.89855e-315 0
0
9 Inverter~
13 330 547 0 2 22
0 27 19
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
4597 0 0
2
5.89855e-315 0
0
9 Inverter~
13 330 511 0 2 22
0 28 20
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
3835 0 0
2
5.89855e-315 0
0
9 Inverter~
13 329 474 0 2 22
0 29 21
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3670 0 0
2
5.89855e-315 0
0
8 Hex Key~
166 141 308 0 11 12
0 32 33 34 35 0 0 0 0 0
9 57
0
0 0 4640 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
5616 0 0
2
5.89855e-315 0
0
8 Hex Key~
166 137 84 0 11 12
0 36 37 38 39 0 0 0 0 0
0 48
0
0 0 4640 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
9323 0 0
2
5.89855e-315 0
0
6 74LS83
105 245 392 0 14 29
0 35 34 33 32 30 30 31 31 30
29 28 27 26 41
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U2
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
317 0 0
2
5.89855e-315 0
0
6 74LS83
105 245 193 0 14 29
0 39 38 37 36 30 30 31 31 30
25 24 23 22 42
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
3108 0 0
2
5.89855e-315 0
0
53
13 1 2 0 0 8320 0 11 5 0 0 3
709 286
798 286
798 151
12 2 3 0 0 8320 0 11 5 0 0 3
709 277
792 277
792 151
11 3 4 0 0 8320 0 11 5 0 0 3
709 268
786 268
786 151
10 4 5 0 0 8320 0 11 5 0 0 3
709 259
780 259
780 151
1 4 6 0 0 8192 0 1 11 0 0 4
597 233
622 233
622 259
645 259
1 3 6 0 0 4096 0 1 11 0 0 4
597 233
627 233
627 250
645 250
1 2 6 0 0 4096 0 1 11 0 0 4
597 233
632 233
632 241
645 241
1 1 6 0 0 4224 0 1 11 0 0 4
597 233
637 233
637 232
645 232
14 9 7 0 0 4224 0 12 11 0 0 4
506 319
617 319
617 313
645 313
3 8 8 0 0 8320 0 7 11 0 0 4
616 527
622 527
622 295
645 295
3 7 9 0 0 8320 0 8 11 0 0 4
615 474
627 474
627 286
645 286
3 6 10 0 0 8320 0 9 11 0 0 4
613 421
632 421
632 277
645 277
3 5 11 0 0 8320 0 10 11 0 0 4
612 367
637 367
637 268
645 268
2 2 12 0 0 8320 0 6 7 0 0 4
533 370
539 370
539 536
567 536
2 2 12 0 0 0 0 6 8 0 0 4
533 370
548 370
548 483
566 483
2 2 12 0 0 0 0 6 9 0 0 4
533 370
541 370
541 430
564 430
2 2 12 0 0 0 0 6 10 0 0 4
533 370
555 370
555 376
563 376
14 1 7 0 0 0 0 12 6 0 0 6
506 319
510 319
510 356
492 356
492 370
497 370
13 1 13 0 0 8320 0 12 7 0 0 4
506 292
544 292
544 518
567 518
12 1 14 0 0 8320 0 12 8 0 0 4
506 283
558 283
558 465
566 465
11 1 15 0 0 8320 0 12 9 0 0 4
506 274
551 274
551 412
564 412
10 1 16 0 0 8320 0 12 10 0 0 4
506 265
555 265
555 358
563 358
1 9 17 0 0 4224 0 2 12 0 0 4
356 287
414 287
414 319
442 319
2 8 18 0 0 8320 0 13 12 0 0 4
351 584
419 584
419 301
442 301
2 7 19 0 0 8320 0 14 12 0 0 4
351 547
424 547
424 292
442 292
2 6 20 0 0 8320 0 15 12 0 0 4
351 511
429 511
429 283
442 283
2 5 21 0 0 8320 0 16 12 0 0 4
350 474
434 474
434 274
442 274
13 4 22 0 0 4224 0 20 12 0 0 4
277 211
419 211
419 265
442 265
12 3 23 0 0 4224 0 20 12 0 0 4
277 202
424 202
424 256
442 256
11 2 24 0 0 4224 0 20 12 0 0 4
277 193
429 193
429 247
442 247
10 1 25 0 0 4224 0 20 12 0 0 4
277 184
434 184
434 238
442 238
13 1 26 0 0 8320 0 19 13 0 0 4
277 410
292 410
292 584
315 584
12 1 27 0 0 8320 0 19 14 0 0 4
277 401
297 401
297 547
315 547
11 1 28 0 0 8320 0 19 15 0 0 4
277 392
302 392
302 511
315 511
10 1 29 0 0 8320 0 19 16 0 0 4
277 383
306 383
306 474
314 474
1 5 30 0 0 8320 0 3 20 0 0 4
155 427
170 427
170 193
213 193
1 6 30 0 0 0 0 3 20 0 0 4
155 427
175 427
175 202
213 202
1 5 30 0 0 0 0 3 19 0 0 4
155 427
180 427
180 392
213 392
1 6 30 0 0 0 0 3 19 0 0 4
155 427
185 427
185 401
213 401
1 9 30 0 0 0 0 3 20 0 0 4
155 427
200 427
200 238
213 238
1 9 30 0 0 0 0 3 19 0 0 4
155 427
205 427
205 437
213 437
1 8 31 0 0 8320 0 4 19 0 0 4
151 228
190 228
190 419
213 419
1 7 31 0 0 0 0 4 19 0 0 4
151 228
195 228
195 410
213 410
1 8 31 0 0 0 0 4 20 0 0 4
151 228
200 228
200 220
213 220
1 7 31 0 0 0 0 4 20 0 0 4
151 228
205 228
205 211
213 211
1 4 32 0 0 8320 0 17 19 0 0 3
150 332
150 383
213 383
2 3 33 0 0 8320 0 17 19 0 0 3
144 332
144 374
213 374
3 2 34 0 0 8320 0 17 19 0 0 3
138 332
138 365
213 365
4 1 35 0 0 8320 0 17 19 0 0 3
132 332
132 356
213 356
1 4 36 0 0 4224 0 18 20 0 0 3
146 108
146 184
213 184
2 3 37 0 0 8320 0 18 20 0 0 3
140 108
140 175
213 175
3 2 38 0 0 8320 0 18 20 0 0 3
134 108
134 166
213 166
4 1 39 0 0 8320 0 18 20 0 0 3
128 108
128 157
213 157
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
407 81 596 105
417 89 585 105
21 XS-3 SUBTRACTOR (1'S)
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
