CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
30
13 Logic Switch~
5 79 501 0 1 11
0 5
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 80 431 0 1 11
0 7
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 82 356 0 1 11
0 6
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 88 200 0 1 11
0 18
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 87 140 0 1 11
0 20
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 87 74 0 1 11
0 19
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
5.89855e-315 0
0
5 4073~
219 412 493 0 4 22
0 4 3 2 28
0
0 0 608 0
4 4073
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 512 3 2 2 0
1 U
8901 0 0
2
5.89855e-315 0
0
5 4082~
219 411 357 0 5 22
0 11 10 9 8 29
0
0 0 608 0
4 4082
-7 -24 21 -16
4 U10A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 512 2 1 10 0
1 U
7361 0 0
2
5.89855e-315 0
0
5 4071~
219 304 520 0 3 22
0 6 5 2
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U8C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 8 0
1 U
4747 0 0
2
5.89855e-315 0
0
5 4071~
219 304 454 0 3 22
0 7 5 3
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U8B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 8 0
1 U
972 0 0
2
5.89855e-315 0
0
5 4071~
219 302 386 0 3 22
0 6 7 4
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U8A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 8 0
1 U
3472 0 0
2
5.89855e-315 0
0
9 Inverter~
13 144 482 0 2 22
0 5 12
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U3F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 3 0
1 U
9998 0 0
2
5.89855e-315 0
0
9 Inverter~
13 145 413 0 2 22
0 7 14
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U3E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 3 0
1 U
3536 0 0
2
5.89855e-315 0
0
9 Inverter~
13 146 336 0 2 22
0 6 13
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U3D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 3 0
1 U
4597 0 0
2
5.89855e-315 0
0
8 3-In OR~
219 211 540 0 4 22
0 13 12 7 8
0
0 0 608 0
4 4075
-14 -24 14 -16
3 U7B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 7 0
1 U
3835 0 0
2
5.89855e-315 0
0
8 3-In OR~
219 213 484 0 4 22
0 13 14 5 9
0
0 0 608 0
4 4075
-14 -24 14 -16
3 U7A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 7 0
1 U
3670 0 0
2
5.89855e-315 0
0
8 3-In OR~
219 213 425 0 4 22
0 6 14 12 10
0
0 0 608 0
4 4075
-14 -24 14 -16
3 U5C
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 5 0
1 U
5616 0 0
2
5.89855e-315 0
0
8 3-In OR~
219 213 360 0 4 22
0 6 7 5 11
0
0 0 608 0
4 4075
-14 -24 14 -16
3 U5B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 5 0
1 U
9323 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 316 219 0 3 22
0 19 18 17
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U6C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
317 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 314 146 0 3 22
0 20 18 16
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U6B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
3108 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 312 74 0 3 22
0 19 20 15
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
4299 0 0
2
5.89855e-315 0
0
8 3-In OR~
219 387 200 0 4 22
0 15 16 17 30
0
0 0 608 0
4 4075
-14 -24 14 -16
3 U5A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 512 3 1 5 0
1 U
9672 0 0
2
5.89855e-315 0
0
8 4-In OR~
219 391 66 0 5 22
0 24 23 22 21 31
0
0 0 608 0
4 4072
-14 -24 14 -16
3 U4A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 512 2 1 4 0
1 U
7876 0 0
2
5.89855e-315 0
0
9 Inverter~
13 142 182 0 2 22
0 18 25
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U3C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
6369 0 0
2
5.89855e-315 0
0
9 Inverter~
13 141 121 0 2 22
0 20 26
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U3B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
9172 0 0
2
5.89855e-315 0
0
9 Inverter~
13 142 55 0 2 22
0 19 27
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
7100 0 0
2
5.89855e-315 0
0
5 4073~
219 227 248 0 4 22
0 19 26 25 21
0
0 0 608 0
4 4073
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 2 0
1 U
3820 0 0
2
5.89855e-315 0
0
5 4073~
219 230 178 0 4 22
0 27 26 18 22
0
0 0 608 0
4 4073
-7 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 1 0
1 U
7678 0 0
2
5.89855e-315 0
0
5 4073~
219 230 109 0 4 22
0 27 20 25 23
0
0 0 608 0
4 4073
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 1 0
1 U
961 0 0
2
5.89855e-315 0
0
5 4073~
219 232 42 0 4 22
0 19 20 18 24
0
0 0 608 0
4 4073
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 1 0
1 U
3178 0 0
2
5.89855e-315 0
0
56
3 3 2 0 0 4224 0 9 7 0 0 4
337 520
380 520
380 502
388 502
3 2 3 0 0 8320 0 10 7 0 0 4
337 454
375 454
375 493
388 493
3 1 4 0 0 8320 0 11 7 0 0 4
335 386
365 386
365 484
388 484
1 2 5 0 0 12288 0 1 9 0 0 6
91 501
184 501
184 560
283 560
283 529
291 529
1 1 6 0 0 8320 0 3 9 0 0 4
94 356
171 356
171 511
291 511
1 2 5 0 0 4096 0 1 10 0 0 4
91 501
196 501
196 463
291 463
1 1 7 0 0 12288 0 2 10 0 0 4
92 431
181 431
181 445
291 445
1 2 7 0 0 0 0 2 11 0 0 4
92 431
196 431
196 395
289 395
1 1 6 0 0 0 0 3 11 0 0 6
94 356
196 356
196 380
281 380
281 377
289 377
4 4 8 0 0 8320 0 15 8 0 0 4
244 540
369 540
369 371
387 371
4 3 9 0 0 4224 0 16 8 0 0 4
246 484
379 484
379 362
387 362
4 2 10 0 0 4224 0 17 8 0 0 4
246 425
374 425
374 353
387 353
4 1 11 0 0 4224 0 18 8 0 0 4
246 360
379 360
379 344
387 344
1 3 7 0 0 8320 0 2 15 0 0 4
92 431
170 431
170 549
198 549
2 2 12 0 0 8320 0 12 15 0 0 4
165 482
180 482
180 540
199 540
2 1 13 0 0 8320 0 14 15 0 0 4
167 336
175 336
175 531
198 531
1 3 5 0 0 0 0 1 16 0 0 4
91 501
192 501
192 493
200 493
2 2 14 0 0 8320 0 13 16 0 0 4
166 413
172 413
172 484
201 484
2 1 13 0 0 0 0 14 16 0 0 4
167 336
172 336
172 475
200 475
2 3 12 0 0 0 0 12 17 0 0 4
165 482
192 482
192 434
200 434
2 2 14 0 0 0 0 13 17 0 0 4
166 413
177 413
177 425
201 425
1 1 6 0 0 0 0 3 17 0 0 4
94 356
182 356
182 416
200 416
1 1 5 0 0 0 0 1 12 0 0 4
91 501
121 501
121 482
129 482
1 1 7 0 0 0 0 2 13 0 0 4
92 431
122 431
122 413
130 413
1 1 6 0 0 0 0 3 14 0 0 4
94 356
123 356
123 336
131 336
1 3 5 0 0 8320 0 1 18 0 0 4
91 501
187 501
187 369
200 369
1 2 7 0 0 0 0 2 18 0 0 4
92 431
192 431
192 360
201 360
1 1 6 0 0 0 0 3 18 0 0 4
94 356
192 356
192 351
200 351
3 1 15 0 0 8320 0 21 22 0 0 4
333 74
351 74
351 191
374 191
3 2 16 0 0 8320 0 20 22 0 0 4
335 146
366 146
366 200
375 200
3 3 17 0 0 4224 0 19 22 0 0 4
337 219
366 219
366 209
374 209
1 2 18 0 0 4096 0 4 19 0 0 4
100 200
279 200
279 228
292 228
1 1 19 0 0 4096 0 6 19 0 0 4
99 74
274 74
274 210
292 210
1 2 18 0 0 4224 0 4 20 0 0 4
100 200
282 200
282 155
290 155
1 1 20 0 0 4096 0 5 20 0 0 4
99 140
277 140
277 137
290 137
1 2 20 0 0 4224 0 5 21 0 0 4
99 140
280 140
280 83
288 83
1 1 19 0 0 4224 0 6 21 0 0 4
99 74
280 74
280 65
288 65
4 4 21 0 0 8320 0 27 23 0 0 4
248 248
356 248
356 80
374 80
4 3 22 0 0 4224 0 28 23 0 0 4
251 178
361 178
361 71
374 71
4 2 23 0 0 4224 0 29 23 0 0 4
251 109
366 109
366 62
374 62
4 1 24 0 0 4224 0 30 23 0 0 4
253 42
366 42
366 53
374 53
2 3 25 0 0 8320 0 24 27 0 0 4
163 182
195 182
195 257
203 257
2 2 26 0 0 8320 0 25 27 0 0 4
162 121
170 121
170 248
203 248
1 1 19 0 0 0 0 6 27 0 0 4
99 74
170 74
170 239
203 239
1 3 18 0 0 0 0 4 28 0 0 4
100 200
198 200
198 187
206 187
2 2 26 0 0 0 0 25 28 0 0 4
162 121
173 121
173 178
206 178
2 1 27 0 0 8320 0 26 28 0 0 4
163 55
178 55
178 169
206 169
2 3 25 0 0 0 0 24 29 0 0 4
163 182
183 182
183 118
206 118
1 2 20 0 0 0 0 5 29 0 0 4
99 140
198 140
198 109
206 109
2 1 27 0 0 0 0 26 29 0 0 4
163 55
183 55
183 100
206 100
1 1 18 0 0 0 0 4 24 0 0 4
100 200
119 200
119 182
127 182
1 1 20 0 0 0 0 5 25 0 0 4
99 140
118 140
118 121
126 121
1 1 19 0 0 0 0 6 26 0 0 4
99 74
119 74
119 55
127 55
1 3 18 0 0 0 0 4 30 0 0 4
100 200
190 200
190 51
208 51
1 2 20 0 0 0 0 5 30 0 0 4
99 140
195 140
195 42
208 42
1 1 19 0 0 0 0 6 30 0 0 4
99 74
200 74
200 33
208 33
7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
182 579 283 603
192 587 272 603
10 FULL ADDER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
422 49 467 73
432 57 456 73
3 Sum
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
414 181 475 205
424 189 464 205
5 Carry
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
487 113 572 137
497 121 561 137
8 SOP Form
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
428 341 473 365
438 349 462 365
3 SUM
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
430 477 491 501
440 485 480 501
5 CARRY
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
506 400 591 424
516 408 580 424
8 POS Form
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
