CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
15
13 Logic Switch~
5 71 363 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43335.1 0
0
13 Logic Switch~
5 71 94 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 69 228 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3124 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 70 177 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 72 51 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8157 0 0
2
5.89859e-315 0
0
14 Logic Display~
6 549 482 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5572 0 0
2
43335.1 0
0
14 Logic Display~
6 444 484 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8901 0 0
2
43335.1 0
0
14 Logic Display~
6 321 487 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7361 0 0
2
43335.1 0
0
14 Logic Display~
6 168 490 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4747 0 0
2
43335.1 0
0
9 2-In AND~
219 350 278 0 3 22
0 11 12 5
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1D
-13 -12 8 -4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
972 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 242 277 0 3 22
0 11 13 8
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1C
-12 -11 9 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3472 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 202 277 0 3 22
0 14 12 9
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1B
-12 -11 9 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
9998 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 133 276 0 3 22
0 14 13 10
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1A
-12 -11 9 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3536 0 0
2
5.89859e-315 0
0
2 FA
94 222 352 0 5 11
0 8 9 4 6 7
2 FA
4 0 688 0
0
2 U2
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
4597 0 0
2
43334.9 0
0
2 FA
94 348 351 0 5 11
0 5 6 4 2 3
2 FA
5 0 688 0
0
2 U3
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
3835 0 0
2
43334.9 0
0
22
4 1 2 0 0 8320 0 15 6 0 0 5
381 369
515 369
515 522
549 522
549 500
5 1 3 0 0 8320 0 15 7 0 0 5
381 351
415 351
415 521
444 521
444 502
0 3 4 0 0 8320 0 0 15 7 0 4
114 370
114 395
315 395
315 369
3 1 5 0 0 4224 0 10 15 0 0 4
348 301
295 301
295 351
315 351
4 2 6 0 0 4224 0 14 15 0 0 4
255 370
307 370
307 360
315 360
5 1 7 0 0 8320 0 14 8 0 0 5
255 352
284 352
284 521
321 521
321 505
1 3 4 0 0 16 0 1 14 0 0 3
83 363
83 370
189 370
3 1 8 0 0 8320 0 11 14 0 0 5
240 300
240 311
174 311
174 352
189 352
3 2 9 0 0 8320 0 12 14 0 0 4
200 300
162 300
162 361
189 361
3 1 10 0 0 4224 0 13 9 0 0 4
131 299
131 521
168 521
168 508
1 0 11 0 0 4096 0 10 0 0 20 2
357 256
357 177
2 0 12 0 0 4096 0 10 0 0 22 2
339 256
339 51
1 0 11 0 0 0 0 11 0 0 20 2
249 255
249 177
2 0 13 0 0 4096 0 11 0 0 21 2
231 255
231 94
1 0 14 0 0 4096 0 12 0 0 19 2
209 255
209 228
2 0 12 0 0 0 0 12 0 0 22 2
191 255
191 51
1 0 14 0 0 0 0 13 0 0 19 2
140 254
140 228
2 0 13 0 0 0 0 13 0 0 21 2
122 254
122 94
1 0 14 0 0 4224 0 3 0 0 0 2
81 228
523 228
1 0 11 0 0 4224 0 4 0 0 0 2
82 177
523 177
1 0 13 0 0 4224 0 2 0 0 0 2
83 94
524 94
1 0 12 0 0 4224 0 5 0 0 0 2
84 51
524 51
8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
533 530 570 554
543 538 559 554
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
426 528 463 552
436 536 452 552
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
303 530 340 554
313 538 329 554
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
150 533 187 557
160 541 176 557
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
18 32 55 56
28 40 44 56
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
16 75 53 99
26 83 42 99
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
15 156 52 180
25 164 41 180
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
14 204 51 228
24 212 40 228
2 B0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
