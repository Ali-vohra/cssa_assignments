CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
180 70 30 160 10
176 80 1534 843
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
17
13 Logic Switch~
5 536 191 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43319.7 0
0
13 Logic Switch~
5 332 301 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89855e-315 5.26354e-315
0
9 Inverter~
13 462 362 0 2 22
0 3 8
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
3124 0 0
2
43319.7 0
0
5 4030~
219 536 497 0 3 22
0 9 8 4
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U4D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 2 0
1 U
3421 0 0
2
43319.7 0
0
5 4030~
219 539 445 0 3 22
0 10 8 5
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U4C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
8157 0 0
2
43319.7 1
0
5 4030~
219 541 394 0 3 22
0 11 8 6
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U4B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
5572 0 0
2
43319.7 0
0
5 4030~
219 539 341 0 3 22
0 12 8 7
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U4A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
8901 0 0
2
43319.7 0
0
14 Logic Display~
6 968 297 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7361 0 0
2
5.89855e-315 5.30499e-315
0
12 Hex Display~
7 861 160 0 18 19
10 14 15 16 17 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
4747 0 0
2
5.89855e-315 5.32571e-315
0
6 74LS83
105 643 270 0 14 29
0 7 6 5 4 2 2 2 2 3
17 16 15 14 13
0
0 0 4848 0
7 74LS83A
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
972 0 0
2
5.89855e-315 5.34643e-315
0
5 4049~
219 265 449 0 2 22
0 20 19
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 1 0
1 U
3472 0 0
2
5.89855e-315 5.3568e-315
0
5 4049~
219 265 410 0 2 22
0 22 21
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 1 0
1 U
9998 0 0
2
5.89855e-315 5.36716e-315
0
5 4049~
219 267 371 0 2 22
0 24 23
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 1 0
1 U
3536 0 0
2
5.89855e-315 5.37752e-315
0
5 4049~
219 267 333 0 2 22
0 26 25
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 1 0
1 U
4597 0 0
2
5.89855e-315 5.38788e-315
0
8 Hex Key~
166 205 170 0 11 12
0 20 22 24 26 0 0 0 0 0
3 51
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3835 0 0
2
5.89855e-315 5.39306e-315
0
8 Hex Key~
166 310 171 0 11 12
0 27 28 29 30 0 0 0 0 0
2 50
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3670 0 0
2
5.89855e-315 5.39824e-315
0
6 74LS83
105 451 273 0 14 29
0 30 29 28 27 25 23 21 19 18
12 11 10 9 3
0
0 0 4848 0
7 74LS83A
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
5616 0 0
2
5.89855e-315 5.40342e-315
0
36
8 1 2 0 0 8320 0 10 1 0 0 4
611 297
562 297
562 191
548 191
1 7 2 0 0 0 0 1 10 0 0 4
548 191
593 191
593 288
611 288
6 1 2 0 0 0 0 10 1 0 0 4
611 279
557 279
557 191
548 191
1 5 2 0 0 0 0 1 10 0 0 4
548 191
598 191
598 270
611 270
14 9 3 0 0 4224 0 17 10 0 0 4
483 318
598 318
598 315
611 315
4 3 4 0 0 8320 0 10 4 0 0 4
611 261
579 261
579 497
569 497
3 3 5 0 0 8320 0 10 5 0 0 4
611 252
585 252
585 445
572 445
2 3 6 0 0 8320 0 10 6 0 0 4
611 243
582 243
582 394
574 394
3 1 7 0 0 8320 0 7 10 0 0 4
572 341
603 341
603 234
611 234
2 2 8 0 0 8320 0 3 4 0 0 4
483 362
487 362
487 506
520 506
2 2 8 0 0 0 0 3 5 0 0 4
483 362
490 362
490 454
523 454
2 2 8 0 0 0 0 3 6 0 0 4
483 362
497 362
497 403
525 403
2 2 8 0 0 0 0 3 7 0 0 4
483 362
515 362
515 350
523 350
14 1 3 0 0 0 0 17 3 0 0 6
483 318
487 318
487 377
439 377
439 362
447 362
13 1 9 0 0 8320 0 17 4 0 0 4
483 291
502 291
502 488
520 488
12 1 10 0 0 8320 0 17 5 0 0 4
483 282
505 282
505 436
523 436
11 1 11 0 0 8320 0 17 6 0 0 4
483 273
512 273
512 385
525 385
10 1 12 0 0 8320 0 17 7 0 0 4
483 264
515 264
515 332
523 332
14 1 13 0 0 4224 0 10 8 0 0 5
675 315
956 315
956 323
968 323
968 315
13 1 14 0 0 4224 0 10 9 0 0 3
675 288
870 288
870 184
12 2 15 0 0 4224 0 10 9 0 0 3
675 279
864 279
864 184
11 3 16 0 0 4224 0 10 9 0 0 3
675 270
858 270
858 184
10 4 17 0 0 4224 0 10 9 0 0 3
675 261
852 261
852 184
1 9 18 0 0 4224 0 2 17 0 0 4
344 301
391 301
391 318
419 318
2 8 19 0 0 8320 0 11 17 0 0 4
286 449
396 449
396 300
419 300
1 1 20 0 0 4224 0 15 11 0 0 3
214 194
214 449
250 449
2 7 21 0 0 8320 0 12 17 0 0 4
286 410
401 410
401 291
419 291
2 1 22 0 0 4224 0 15 12 0 0 3
208 194
208 410
250 410
2 6 23 0 0 4224 0 13 17 0 0 4
288 371
406 371
406 282
419 282
3 1 24 0 0 4224 0 15 13 0 0 3
202 194
202 371
252 371
2 5 25 0 0 4224 0 14 17 0 0 4
288 333
411 333
411 273
419 273
4 1 26 0 0 4224 0 15 14 0 0 3
196 194
196 333
252 333
1 4 27 0 0 8320 0 16 17 0 0 3
319 195
319 264
419 264
2 3 28 0 0 8320 0 16 17 0 0 3
313 195
313 255
419 255
3 2 29 0 0 8320 0 16 17 0 0 3
307 195
307 246
419 246
4 1 30 0 0 8320 0 16 17 0 0 3
301 195
301 237
419 237
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
423 78 620 102
433 86 609 102
22 BINARY SUBTRACTOR(1'S)
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
