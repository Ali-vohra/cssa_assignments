CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
13
13 Logic Switch~
5 391 261 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V3
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7361 0 0
2
43362 0
0
13 Logic Switch~
5 275 262 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V2
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4747 0 0
2
43362 0
0
13 Logic Switch~
5 125 123 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
972 0 0
2
43362 0
0
14 Logic Display~
6 641 183 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3472 0 0
2
43362 0
0
14 Logic Display~
6 642 128 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9998 0 0
2
43362 0
0
14 Logic Display~
6 641 78 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3536 0 0
2
43362 0
0
14 Logic Display~
6 641 25 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4597 0 0
2
43362 0
0
5 4073~
219 485 194 0 4 22
0 10 7 6 2
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 3 0
1 U
3835 0 0
2
43362 0
0
5 4073~
219 486 144 0 4 22
0 10 7 8 3
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 2 0
1 U
3670 0 0
2
43362 0
0
5 4073~
219 487 96 0 4 22
0 10 9 6 4
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 2 0
1 U
5616 0 0
2
43362 0
0
5 4073~
219 488 47 0 4 22
0 10 9 8 5
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 2 0
1 U
9323 0 0
2
43362 0
0
9 Inverter~
13 360 223 0 2 22
0 9 7
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U1B
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
317 0 0
2
43362 0
0
9 Inverter~
13 242 221 0 2 22
0 8 6
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U1A
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3108 0 0
2
43362 0
0
22
4 1 2 0 0 4224 0 8 4 0 0 5
506 194
629 194
629 209
641 209
641 201
4 1 3 0 0 4224 0 9 5 0 0 5
507 144
630 144
630 154
642 154
642 146
4 1 4 0 0 4224 0 10 6 0 0 5
508 96
629 96
629 104
641 104
641 96
4 1 5 0 0 4224 0 11 7 0 0 3
509 47
641 47
641 43
3 2 6 0 0 4096 0 8 13 0 0 2
461 203
245 203
2 0 7 0 0 4096 0 8 0 0 19 2
461 194
363 194
3 0 8 0 0 4096 0 9 0 0 17 2
462 153
276 153
2 0 7 0 0 4096 0 9 0 0 19 2
462 144
363 144
3 0 6 0 0 4224 0 10 0 0 20 2
463 105
245 105
2 0 9 0 0 4096 0 10 0 0 18 2
463 96
392 96
3 0 8 0 0 4096 0 11 0 0 17 2
464 56
276 56
2 0 9 0 0 4096 0 11 0 0 18 2
464 47
392 47
1 1 10 0 0 4096 0 8 3 0 0 4
461 185
161 185
161 123
137 123
1 1 10 0 0 4096 0 9 3 0 0 4
462 135
156 135
156 123
137 123
1 1 10 0 0 4096 0 10 3 0 0 4
463 87
151 87
151 123
137 123
1 1 10 0 0 4224 0 11 3 0 0 4
464 38
146 38
146 123
137 123
1 0 8 0 0 4224 0 2 0 0 0 2
276 249
276 19
1 0 9 0 0 4224 0 1 0 0 0 2
392 248
392 20
2 0 7 0 0 4224 0 12 0 0 0 2
363 205
363 19
2 0 6 0 0 0 0 13 0 0 0 2
245 203
245 18
1 1 9 0 0 0 0 1 12 0 0 4
392 248
392 243
363 243
363 241
1 1 8 0 0 0 0 2 13 0 0 4
276 249
276 241
245 241
245 239
7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
665 169 702 193
675 177 691 193
2 D0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
665 113 702 137
675 121 691 137
2 D1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
663 62 700 86
673 70 689 86
2 D2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
661 9 698 33
671 17 687 33
2 D3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
375 280 412 304
385 288 401 304
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
258 280 295 304
268 288 284 304
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
70 100 107 124
80 108 96 124
2 A0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
