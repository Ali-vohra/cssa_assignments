CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
30 20 30 70 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
27
13 Logic Switch~
5 83 804 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V16
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9323 0 0
2
43355.1 0
0
13 Logic Switch~
5 84 753 0 1 11
0 16
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V15
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
317 0 0
2
43355.1 0
0
13 Logic Switch~
5 84 704 0 1 11
0 17
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V14
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3108 0 0
2
43355.1 0
0
13 Logic Switch~
5 86 659 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V13
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4299 0 0
2
43355.1 0
0
13 Logic Switch~
5 86 612 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V12
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9672 0 0
2
43355.1 0
0
13 Logic Switch~
5 88 561 0 1 11
0 20
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V11
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7876 0 0
2
43355.1 0
0
13 Logic Switch~
5 89 512 0 1 11
0 21
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V10
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6369 0 0
2
43355.1 0
0
13 Logic Switch~
5 89 464 0 1 11
0 22
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9172 0 0
2
43355.1 0
0
13 Logic Switch~
5 89 418 0 1 11
0 23
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7100 0 0
2
43355.1 0
0
13 Logic Switch~
5 89 366 0 1 11
0 24
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3820 0 0
2
43355.1 0
0
13 Logic Switch~
5 89 321 0 1 11
0 25
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7678 0 0
2
43355.1 0
0
13 Logic Switch~
5 87 269 0 1 11
0 26
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
961 0 0
2
43355.1 0
0
13 Logic Switch~
5 87 214 0 1 11
0 27
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3178 0 0
2
43355.1 0
0
13 Logic Switch~
5 85 160 0 1 11
0 28
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3409 0 0
2
43355.1 0
0
13 Logic Switch~
5 85 107 0 1 11
0 29
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3951 0 0
2
43355.1 0
0
13 Logic Switch~
5 85 54 0 10 11
0 30 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8885 0 0
2
43355.1 0
0
14 Logic Display~
6 842 353 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3780 0 0
2
43355.1 0
0
14 Logic Display~
6 842 293 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9265 0 0
2
43355.1 0
0
14 Logic Display~
6 841 235 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9442 0 0
2
43355.1 0
0
14 Logic Display~
6 841 178 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9424 0 0
2
43355.1 0
0
8 2-In OR~
219 587 396 0 3 22
0 7 6 2
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
9968 0 0
2
43355.1 0
0
8 2-In OR~
219 589 346 0 3 22
0 9 8 3
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
9281 0 0
2
43355.1 0
0
8 2-In OR~
219 591 291 0 3 22
0 11 10 4
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
8464 0 0
2
43355.1 0
0
9 2-In AND~
219 598 242 0 3 22
0 13 12 5
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
7168 0 0
2
43355.1 0
0
9 Inverter~
13 476 482 0 2 22
0 14 12
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3171 0 0
2
43355.1 0
0
8 8-3 ENC~
94 413 151 0 12 25
0 30 29 28 27 26 25 24 23 13
7 9 11
7 8-3 ENC
1 0 560 0
0
2 U1
-3 -77 11 -69
0
0
0
0
0
0
25

0 1 2 3 4 5 6 7 8 9
12 13 14 1 2 3 4 5 6 7
8 9 12 13 14 0
0 0 0 0 0 0 0 0
1 U
4139 0 0
2
43355.1 0
0
8 8-3 ENC~
94 412 428 0 12 25
0 22 21 20 19 18 17 16 15 14
6 8 10
7 8-3 ENC
2 0 560 0
0
2 U2
-3 -77 11 -69
0
0
0
0
0
0
25

0 1 2 3 4 5 6 7 8 9
12 13 14 1 2 3 4 5 6 7
8 9 12 13 14 0
0 0 0 0 0 0 0 0
1 U
6435 0 0
2
43355.1 0
0
29
3 1 2 0 0 4224 0 21 17 0 0 3
620 396
842 396
842 371
3 1 3 0 0 4224 0 22 18 0 0 5
622 346
830 346
830 319
842 319
842 311
3 1 4 0 0 4224 0 23 19 0 0 5
624 291
830 291
830 261
841 261
841 253
3 1 5 0 0 4224 0 24 20 0 0 5
619 242
829 242
829 204
841 204
841 196
10 2 6 0 0 4224 0 27 21 0 0 4
462 441
556 441
556 405
574 405
10 1 7 0 0 8320 0 26 21 0 0 4
463 164
556 164
556 387
574 387
11 2 8 0 0 4224 0 27 22 0 0 4
462 428
563 428
563 355
576 355
11 1 9 0 0 8320 0 26 22 0 0 4
463 151
563 151
563 337
576 337
12 2 10 0 0 8320 0 27 23 0 0 4
462 415
570 415
570 300
578 300
12 1 11 0 0 8320 0 26 23 0 0 4
463 138
570 138
570 282
578 282
2 2 12 0 0 8320 0 25 24 0 0 4
497 482
566 482
566 251
574 251
9 1 13 0 0 4224 0 26 24 0 0 4
463 205
566 205
566 233
574 233
1 9 14 0 0 4224 0 25 27 0 0 2
461 482
462 482
1 8 15 0 0 8320 0 1 27 0 0 4
95 804
332 804
332 482
370 482
1 7 16 0 0 8320 0 2 27 0 0 4
96 753
362 753
362 468
370 468
1 6 17 0 0 8320 0 3 27 0 0 4
96 704
337 704
337 455
370 455
1 5 18 0 0 4224 0 4 27 0 0 4
98 659
342 659
342 441
370 441
1 4 19 0 0 4224 0 5 27 0 0 4
98 612
347 612
347 428
370 428
1 3 20 0 0 4224 0 6 27 0 0 4
100 561
352 561
352 415
370 415
1 2 21 0 0 4224 0 7 27 0 0 4
101 512
357 512
357 401
370 401
1 1 22 0 0 4224 0 8 27 0 0 4
101 464
362 464
362 388
370 388
1 8 23 0 0 4224 0 9 26 0 0 4
101 418
343 418
343 205
371 205
1 7 24 0 0 4224 0 10 26 0 0 4
101 366
348 366
348 191
371 191
1 6 25 0 0 4224 0 11 26 0 0 4
101 321
353 321
353 178
371 178
1 5 26 0 0 4224 0 12 26 0 0 4
99 269
363 269
363 164
371 164
1 4 27 0 0 4224 0 13 26 0 0 4
99 214
358 214
358 151
371 151
1 3 28 0 0 4224 0 14 26 0 0 4
97 160
363 160
363 138
371 138
1 2 29 0 0 4224 0 15 26 0 0 4
97 107
358 107
358 124
371 124
1 1 30 0 0 4224 0 16 26 0 0 4
97 54
363 54
363 111
371 111
20
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
863 342 890 366
868 346 884 362
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
862 281 889 305
867 285 883 301
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
863 224 890 248
868 228 884 244
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
863 167 890 191
868 171 884 187
2 A3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
38 787 65 811
43 791 59 807
2 D0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
37 737 64 761
42 741 58 757
2 D1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
38 688 65 712
43 692 59 708
2 D2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
38 643 65 667
43 647 59 663
2 D3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
38 597 65 621
43 601 59 617
2 D4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
38 546 65 570
43 550 59 566
2 D5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
38 496 65 520
43 500 59 516
2 D6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
39 446 66 470
44 450 60 466
2 D7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
38 401 65 425
43 405 59 421
2 D8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
38 350 65 374
43 354 59 370
2 D9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
36 304 71 328
41 308 65 324
3 D10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
34 253 69 277
39 257 63 273
3 D11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
34 197 69 221
39 201 63 217
3 D12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
33 142 68 166
38 146 62 162
3 D13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
32 91 67 115
37 95 61 111
3 D14
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
32 36 67 60
37 40 61 56
3 D15
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
