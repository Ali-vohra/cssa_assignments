CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
130 50 30 130 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
13
13 Logic Switch~
5 772 240 0 1 11
0 3
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 618 369 0 1 11
0 9
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 162 478 0 1 11
0 14
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 169 237 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
5.89855e-315 0
0
12 Hex Display~
7 891 166 0 18 19
10 4 5 6 7 0 0 0 0 0
0 1 1 1 1 0 0 1 3
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
8157 0 0
2
5.89855e-315 0
0
12 Hex Display~
7 810 168 0 18 19
10 2 3 3 3 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
5572 0 0
2
5.89855e-315 0
0
9 Inverter~
13 572 393 0 2 22
0 2 8
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U5A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
8901 0 0
2
5.89855e-315 0
0
6 74LS83
105 713 314 0 14 29
0 8 8 2 9 13 12 11 10 9
7 6 5 4 32
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U4
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
7361 0 0
2
5.89855e-315 0
0
6 74LS83
105 501 317 0 14 29
0 22 21 20 19 18 17 16 15 14
13 12 11 10 2
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U3
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
4747 0 0
2
5.89855e-315 0
0
8 Hex Key~
166 154 342 0 11 12
0 24 25 26 27 0 0 0 0 0
8 56
0
0 0 4640 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
972 0 0
2
5.89855e-315 0
0
8 Hex Key~
166 150 86 0 11 12
0 28 29 30 31 0 0 0 0 0
5 53
0
0 0 4640 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3472 0 0
2
5.89855e-315 0
0
6 74LS83
105 277 442 0 14 29
0 27 26 25 24 14 14 23 14 14
18 17 16 15 33
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U2
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
9998 0 0
2
5.89855e-315 0
0
6 74LS83
105 273 208 0 14 29
0 31 30 29 28 14 14 23 14 14
22 21 20 19 34
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
3536 0 0
2
5.89855e-315 0
0
45
14 1 2 0 0 12416 0 9 6 0 0 5
533 362
599 362
599 200
819 200
819 192
1 2 3 0 0 8320 0 1 6 0 0 3
784 240
813 240
813 192
1 3 3 0 0 0 0 1 6 0 0 3
784 240
807 240
807 192
1 4 3 0 0 0 0 1 6 0 0 3
784 240
801 240
801 192
13 1 4 0 0 4224 0 8 5 0 0 3
745 332
900 332
900 190
12 2 5 0 0 4224 0 8 5 0 0 3
745 323
894 323
894 190
11 3 6 0 0 4224 0 8 5 0 0 3
745 314
888 314
888 190
10 4 7 0 0 4224 0 8 5 0 0 3
745 305
882 305
882 190
14 3 2 0 0 0 0 9 8 0 0 4
533 362
604 362
604 296
681 296
2 2 8 0 0 8192 0 7 8 0 0 4
593 393
658 393
658 287
681 287
2 1 8 0 0 8320 0 7 8 0 0 4
593 393
663 393
663 278
681 278
14 1 2 0 0 0 0 9 7 0 0 4
533 362
549 362
549 393
557 393
1 4 9 0 0 8320 0 2 8 0 0 4
630 369
668 369
668 305
681 305
1 9 9 0 0 0 0 2 8 0 0 4
630 369
673 369
673 359
681 359
13 8 10 0 0 4224 0 9 8 0 0 4
533 335
673 335
673 341
681 341
12 7 11 0 0 4224 0 9 8 0 0 4
533 326
673 326
673 332
681 332
11 6 12 0 0 4224 0 9 8 0 0 4
533 317
673 317
673 323
681 323
10 5 13 0 0 4224 0 9 8 0 0 4
533 308
673 308
673 314
681 314
1 9 14 0 0 12288 0 3 9 0 0 4
174 478
241 478
241 362
469 362
13 8 15 0 0 4224 0 12 9 0 0 4
309 460
446 460
446 344
469 344
12 7 16 0 0 4224 0 12 9 0 0 4
309 451
451 451
451 335
469 335
11 6 17 0 0 4224 0 12 9 0 0 4
309 442
456 442
456 326
469 326
10 5 18 0 0 4224 0 12 9 0 0 4
309 433
461 433
461 317
469 317
13 4 19 0 0 4224 0 13 9 0 0 4
305 226
446 226
446 308
469 308
12 3 20 0 0 4224 0 13 9 0 0 4
305 217
451 217
451 299
469 299
11 2 21 0 0 4224 0 13 9 0 0 4
305 208
456 208
456 290
469 290
10 1 22 0 0 4224 0 13 9 0 0 4
305 199
461 199
461 281
469 281
1 6 14 0 0 8192 0 3 13 0 0 4
174 478
203 478
203 217
241 217
1 5 14 0 0 8320 0 3 13 0 0 4
174 478
208 478
208 208
241 208
1 8 14 0 0 0 0 3 13 0 0 4
174 478
213 478
213 235
241 235
1 9 14 0 0 0 0 3 13 0 0 4
174 478
218 478
218 253
241 253
1 9 14 0 0 0 0 3 12 0 0 4
174 478
222 478
222 487
245 487
1 8 14 0 0 0 0 3 12 0 0 4
174 478
237 478
237 469
245 469
1 6 14 0 0 0 0 3 12 0 0 4
174 478
227 478
227 451
245 451
1 5 14 0 0 0 0 3 12 0 0 4
174 478
232 478
232 442
245 442
1 7 23 0 0 8320 0 4 12 0 0 4
181 237
237 237
237 460
245 460
1 7 23 0 0 0 0 4 13 0 0 4
181 237
233 237
233 226
241 226
1 4 24 0 0 8320 0 10 12 0 0 3
163 366
163 433
245 433
2 3 25 0 0 8320 0 10 12 0 0 3
157 366
157 424
245 424
3 2 26 0 0 8320 0 10 12 0 0 3
151 366
151 415
245 415
4 1 27 0 0 8320 0 10 12 0 0 3
145 366
145 406
245 406
1 4 28 0 0 4224 0 11 13 0 0 3
159 110
159 199
241 199
2 3 29 0 0 8320 0 11 13 0 0 3
153 110
153 190
241 190
3 2 30 0 0 8320 0 11 13 0 0 3
147 110
147 181
241 181
4 1 31 0 0 8320 0 11 13 0 0 3
141 110
141 172
241 172
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
479 99 580 123
489 107 569 123
10 XS-2 ADDER
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
