CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 50 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
60
13 Logic Switch~
5 60 401 0 10 11
0 60 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43334.8 0
0
13 Logic Switch~
5 60 351 0 10 11
0 43 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
43334.8 0
0
13 Logic Switch~
5 60 302 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
43334.8 0
0
13 Logic Switch~
5 60 254 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3421 0 0
2
43334.8 0
0
13 Logic Switch~
5 57 167 0 10 11
0 59 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8157 0 0
2
43334.8 0
0
13 Logic Switch~
5 57 121 0 10 11
0 42 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5572 0 0
2
43334.8 0
0
13 Logic Switch~
5 57 73 0 10 11
0 25 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8901 0 0
2
43334.8 0
0
13 Logic Switch~
5 58 32 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7361 0 0
2
43334.8 0
0
14 Logic Display~
6 1490 1114 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4747 0 0
2
43334.9 0
0
14 Logic Display~
6 1384 1116 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
972 0 0
2
43334.9 0
0
14 Logic Display~
6 1173 1117 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3472 0 0
2
43334.9 0
0
14 Logic Display~
6 944 1120 0 1 2
10 31
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9998 0 0
2
43334.9 0
0
14 Logic Display~
6 687 1120 0 1 2
10 48
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3536 0 0
2
43334.9 0
0
14 Logic Display~
6 418 1118 0 1 2
10 61
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4597 0 0
2
43334.9 0
0
14 Logic Display~
6 287 1121 0 1 2
10 70
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3835 0 0
2
43334.9 0
0
14 Logic Display~
6 149 1122 0 1 2
10 73
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3670 0 0
2
43334.9 0
0
8 2-In OR~
219 1406 545 0 3 22
0 4 3 2
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U20D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
5616 0 0
2
43334.9 0
0
9 2-In AND~
219 1302 444 0 3 22
0 5 6 8
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U14D
-14 -10 14 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
9323 0 0
2
43334.9 0
0
8 2-In OR~
219 1196 714 0 3 22
0 13 12 10
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U20C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
317 0 0
2
43334.9 0
0
8 2-In OR~
219 1196 552 0 3 22
0 15 14 11
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U20B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
3108 0 0
2
43334.9 0
0
9 2-In AND~
219 1125 445 0 3 22
0 6 25 19
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U14C
-15 -11 13 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
4299 0 0
2
43334.9 0
0
9 2-In AND~
219 1083 446 0 3 22
0 26 5 20
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U14B
-15 -10 13 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
9672 0 0
2
43334.9 0
0
8 2-In OR~
219 968 716 0 3 22
0 28 27 23
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U20A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
7876 0 0
2
43334.9 0
0
8 2-In OR~
219 970 558 0 3 22
0 30 29 24
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
6369 0 0
2
43334.9 0
0
9 2-In AND~
219 907 445 0 3 22
0 6 42 34
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U14A
-15 -10 13 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
9172 0 0
2
43334.9 0
0
9 2-In AND~
219 866 446 0 3 22
0 26 25 36
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U8D
-12 -10 9 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
7100 0 0
2
43334.9 0
0
9 2-In AND~
219 826 446 0 3 22
0 43 5 37
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U8C
-12 -9 9 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
3820 0 0
2
43334.9 0
0
8 2-In OR~
219 703 713 0 3 22
0 45 44 40
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
7678 0 0
2
43334.9 0
0
8 2-In OR~
219 705 561 0 3 22
0 47 46 41
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
961 0 0
2
43334.9 0
0
9 2-In AND~
219 654 447 0 3 22
0 6 59 52
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U8B
-12 -9 9 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3178 0 0
2
43334.9 0
0
9 2-In AND~
219 614 447 0 3 22
0 26 42 53
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U8A
-12 -9 9 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3409 0 0
2
43334.9 0
0
9 2-In AND~
219 572 448 0 3 22
0 43 25 54
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3D
-11 -9 10 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
3951 0 0
2
43334.9 0
0
9 2-In AND~
219 530 449 0 3 22
0 60 5 55
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3C
-11 -8 10 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
8885 0 0
2
43334.9 0
0
8 2-In OR~
219 426 644 0 3 22
0 63 62 57
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3780 0 0
2
43334.8 0
0
9 2-In AND~
219 366 450 0 3 22
0 26 59 66
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3B
-12 -9 9 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
9265 0 0
2
43334.8 0
0
9 2-In AND~
219 320 451 0 3 22
0 43 42 68
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3A
-12 -9 9 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
9442 0 0
2
43334.8 0
0
9 2-In AND~
219 275 451 0 3 22
0 60 25 69
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1D
-12 -8 9 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
9424 0 0
2
43334.8 0
0
9 2-In AND~
219 207 450 0 3 22
0 43 59 71
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1C
-12 -6 9 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
9968 0 0
2
43334.8 0
0
9 2-In AND~
219 158 451 0 3 22
0 60 42 72
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1B
-12 -6 9 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
9281 0 0
2
43334.8 0
0
9 2-In AND~
219 108 450 0 3 22
0 60 59 73
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1A
-12 -5 9 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
8464 0 0
2
43334.8 0
0
2 HA
94 183 532 0 4 9
0 72 71 64 70
2 HA
1 0 656 0
0
2 U2
-7 -28 7 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 U
7168 0 0
2
43334.7 0
0
2 HA
94 317 532 0 4 9
0 69 68 58 67
2 HA
2 0 656 0
0
2 U4
-7 -28 7 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 U
3171 0 0
2
43334.7 0
0
2 HA
94 317 605 0 4 9
0 67 66 63 65
2 HA
3 0 656 0
0
2 U5
-7 -28 7 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 U
4139 0 0
2
43334.7 0
0
2 HA
94 317 678 0 4 9
0 64 65 62 61
2 HA
4 0 656 0
0
2 U6
-7 -28 7 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 U
6435 0 0
2
43334.7 0
0
2 HA
94 596 522 0 4 9
0 58 57 47 56
2 HA
5 0 656 0
0
2 U9
-7 -28 7 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 U
5283 0 0
2
43334.7 0
0
2 HA
94 596 599 0 4 9
0 55 56 46 50
2 HA
6 0 656 0
0
3 U10
-11 -28 10 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 U
6874 0 0
2
43334.7 0
0
2 HA
94 596 672 0 4 9
0 54 53 45 51
2 HA
7 0 656 0
0
3 U11
-11 -28 10 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 U
5305 0 0
2
43334.7 0
0
2 HA
94 596 752 0 4 9
0 52 51 44 49
2 HA
8 0 656 0
0
3 U12
-11 -28 10 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 U
34 0 0
2
43334.7 0
0
2 HA
94 597 836 0 4 9
0 49 50 38 48
2 HA
9 0 656 0
0
3 U13
-11 -28 10 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 U
969 0 0
2
43334.7 0
0
2 HA
94 869 515 0 4 9
0 41 40 30 39
2 HA
10 0 656 0
0
3 U15
-11 -28 10 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 U
8402 0 0
2
43334.7 0
0
2 HA
94 870 594 0 4 9
0 38 39 29 32
2 HA
11 0 656 0
0
3 U16
-11 -28 10 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 U
3751 0 0
2
43334.7 0
0
2 HA
94 870 671 0 4 9
0 37 36 28 35
2 HA
12 0 656 0
0
3 U17
-11 -28 10 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 U
4292 0 0
2
43334.7 0
0
2 HA
94 870 750 0 4 9
0 35 34 27 33
2 HA
13 0 656 0
0
3 U18
-11 -28 10 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 U
6118 0 0
2
43334.7 0
0
2 HA
94 869 831 0 4 9
0 32 33 21 31
2 HA
14 0 656 0
0
3 U19
-11 -28 10 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 U
34 0 0
2
43334.7 0
0
2 HA
94 1104 513 0 4 9
0 24 23 15 22
2 HA
15 0 656 0
0
3 U21
-11 -28 10 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 U
6357 0 0
2
43334.7 0
0
2 HA
94 1104 586 0 4 9
0 21 22 14 17
2 HA
16 0 656 0
0
3 U22
-11 -28 10 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 U
319 0 0
2
43334.7 0
0
2 HA
94 1105 667 0 4 9
0 20 19 13 18
2 HA
17 0 656 0
0
3 U23
-11 -28 10 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 U
3976 0 0
2
43334.7 0
0
2 HA
94 1104 749 0 4 9
0 17 18 12 16
2 HA
18 0 656 0
0
3 U24
-11 -28 10 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 U
7634 0 0
2
43334.7 0
0
2 HA
94 1309 510 0 4 9
0 11 10 4 9
2 HA
19 0 656 0
0
3 U25
-11 -28 10 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 U
523 0 0
2
43334.7 0
0
2 HA
94 1309 588 0 4 9
0 9 8 3 7
2 HA
20 0 656 0
0
3 U26
-11 -28 10 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 U
6748 0 0
2
43334.7 0
0
104
3 1 2 0 0 8320 0 17 9 0 0 5
1439 545
1465 545
1465 1159
1490 1159
1490 1132
3 2 3 0 0 4224 0 60 17 0 0 4
1342 597
1385 597
1385 554
1393 554
3 1 4 0 0 4224 0 59 17 0 0 4
1342 519
1385 519
1385 536
1393 536
1 0 5 0 0 4096 0 18 0 0 104 2
1309 422
1309 32
2 0 6 0 0 4096 0 18 0 0 100 2
1291 422
1291 254
4 1 7 0 0 8320 0 60 10 0 0 5
1342 588
1363 588
1363 1158
1384 1158
1384 1134
3 2 8 0 0 12416 0 18 60 0 0 5
1300 467
1300 475
1247 475
1247 597
1276 597
4 1 9 0 0 12416 0 59 60 0 0 6
1342 510
1362 510
1362 547
1256 547
1256 588
1276 588
3 2 10 0 0 8320 0 19 59 0 0 4
1229 714
1237 714
1237 519
1276 519
3 1 11 0 0 8320 0 20 59 0 0 3
1229 552
1229 510
1276 510
3 2 12 0 0 4224 0 58 19 0 0 4
1137 758
1175 758
1175 723
1183 723
3 1 13 0 0 4224 0 57 19 0 0 4
1138 676
1175 676
1175 705
1183 705
3 2 14 0 0 4224 0 56 20 0 0 4
1137 595
1175 595
1175 561
1183 561
3 1 15 0 0 4224 0 55 20 0 0 4
1137 522
1175 522
1175 543
1183 543
4 1 16 0 0 8320 0 58 11 0 0 5
1137 749
1152 749
1152 1158
1173 1158
1173 1135
4 1 17 0 0 8320 0 56 58 0 0 6
1137 586
1146 586
1146 706
1036 706
1036 749
1071 749
4 2 18 0 0 12416 0 57 58 0 0 6
1138 667
1151 667
1151 699
1030 699
1030 758
1071 758
3 2 19 0 0 12416 0 21 57 0 0 5
1123 468
1123 472
1043 472
1043 676
1072 676
3 1 20 0 0 12416 0 22 57 0 0 5
1081 469
1081 478
1035 478
1035 667
1072 667
3 1 21 0 0 8320 0 54 56 0 0 4
902 840
1023 840
1023 586
1071 586
4 2 22 0 0 12416 0 55 56 0 0 6
1137 513
1150 513
1150 547
1055 547
1055 595
1071 595
3 2 23 0 0 8336 0 23 55 0 0 4
1001 716
1013 716
1013 522
1071 522
3 1 24 0 0 8320 0 24 55 0 0 3
1003 558
1003 513
1071 513
1 0 6 0 0 4096 0 21 0 0 100 2
1132 423
1132 254
2 0 25 0 0 4096 0 21 0 0 103 2
1114 423
1114 73
1 0 26 0 0 4096 0 22 0 0 99 2
1090 424
1090 302
2 0 5 0 0 4096 0 22 0 0 104 2
1072 424
1072 32
3 2 27 0 0 4224 0 53 23 0 0 4
903 759
947 759
947 725
955 725
3 1 28 0 0 4224 0 52 23 0 0 4
903 680
947 680
947 707
955 707
3 2 29 0 0 4224 0 51 24 0 0 4
903 603
949 603
949 567
957 567
3 1 30 0 0 4224 0 50 24 0 0 4
902 524
949 524
949 549
957 549
4 1 31 0 0 8320 0 54 12 0 0 5
902 831
920 831
920 1158
944 1158
944 1138
4 1 32 0 0 8320 0 51 54 0 0 6
903 594
932 594
932 795
806 795
806 831
836 831
4 2 33 0 0 12416 0 53 54 0 0 6
903 750
926 750
926 788
800 788
800 840
836 840
3 2 34 0 0 12416 0 25 53 0 0 7
905 468
905 480
926 480
926 712
804 712
804 759
837 759
4 1 35 0 0 12416 0 52 53 0 0 6
903 671
921 671
921 708
799 708
799 750
837 750
3 2 36 0 0 12416 0 26 52 0 0 5
864 469
864 480
799 480
799 680
837 680
3 1 37 0 0 4224 0 27 52 0 0 3
824 469
824 671
837 671
3 1 38 0 0 8320 0 49 51 0 0 4
630 845
817 845
817 594
837 594
4 2 39 0 0 12416 0 50 51 0 0 6
902 515
920 515
920 550
808 550
808 603
837 603
3 2 40 0 0 8320 0 28 50 0 0 4
736 713
747 713
747 524
836 524
3 1 41 0 0 8320 0 29 50 0 0 3
738 561
738 515
836 515
1 0 6 0 0 0 0 25 0 0 100 2
914 423
914 254
2 0 42 0 0 4096 0 25 0 0 102 2
896 423
896 121
1 0 26 0 0 0 0 26 0 0 99 2
873 424
873 302
2 0 25 0 0 4096 0 26 0 0 103 2
855 424
855 73
1 0 43 0 0 4096 0 27 0 0 98 2
833 424
833 351
2 0 5 0 0 0 0 27 0 0 104 2
815 424
815 32
3 2 44 0 0 4224 0 48 28 0 0 4
629 761
682 761
682 722
690 722
3 1 45 0 0 4224 0 47 28 0 0 4
629 681
682 681
682 704
690 704
3 2 46 0 0 4224 0 46 29 0 0 4
629 608
684 608
684 570
692 570
3 1 47 0 0 4224 0 45 29 0 0 4
629 531
684 531
684 552
692 552
4 1 48 0 0 8320 0 49 13 0 0 5
630 836
667 836
667 1159
687 1159
687 1138
4 1 49 0 0 12416 0 48 49 0 0 6
629 752
659 752
659 797
530 797
530 836
564 836
4 2 50 0 0 8320 0 46 49 0 0 6
629 599
668 599
668 787
520 787
520 845
564 845
4 2 51 0 0 12416 0 47 48 0 0 6
629 672
643 672
643 706
544 706
544 761
563 761
3 1 52 0 0 4224 0 30 48 0 0 5
652 470
652 713
538 713
538 752
563 752
3 2 53 0 0 12416 0 31 47 0 0 5
612 470
612 477
479 477
479 681
563 681
3 1 54 0 0 12416 0 32 47 0 0 5
570 471
570 487
487 487
487 672
563 672
3 1 55 0 0 4224 0 33 46 0 0 3
528 472
528 599
563 599
4 2 56 0 0 12416 0 45 46 0 0 6
629 522
667 522
667 557
543 557
543 608
563 608
3 2 57 0 0 8320 0 34 45 0 0 4
459 644
513 644
513 531
563 531
3 1 58 0 0 4224 0 42 45 0 0 4
350 541
459 541
459 522
563 522
1 0 6 0 0 4096 0 30 0 0 100 2
661 425
661 254
2 0 59 0 0 4096 0 30 0 0 101 2
643 425
643 167
1 0 26 0 0 4096 0 31 0 0 99 2
621 425
621 302
2 0 42 0 0 4096 0 31 0 0 102 2
603 425
603 121
1 0 43 0 0 4096 0 32 0 0 98 2
579 426
579 351
2 0 25 0 0 4096 0 32 0 0 103 2
561 426
561 73
1 0 60 0 0 4096 0 33 0 0 97 2
537 427
537 401
2 0 5 0 0 4096 0 33 0 0 104 2
519 427
519 32
4 1 61 0 0 8320 0 44 14 0 0 5
350 678
380 678
380 1158
418 1158
418 1136
3 2 62 0 0 4224 0 44 34 0 0 4
350 687
405 687
405 653
413 653
3 1 63 0 0 4224 0 43 34 0 0 4
350 614
405 614
405 635
413 635
3 1 64 0 0 8320 0 41 44 0 0 4
216 541
245 541
245 678
284 678
4 2 65 0 0 12416 0 43 44 0 0 6
350 605
379 605
379 640
256 640
256 687
284 687
3 2 66 0 0 4224 0 35 43 0 0 5
364 473
364 572
272 572
272 614
284 614
4 1 67 0 0 12416 0 42 43 0 0 6
350 532
379 532
379 566
257 566
257 605
284 605
3 2 68 0 0 8320 0 36 42 0 0 5
318 474
318 498
258 498
258 541
284 541
3 1 69 0 0 4224 0 37 42 0 0 3
273 474
273 532
284 532
1 0 26 0 0 4096 0 35 0 0 99 2
373 428
373 302
2 0 59 0 0 4096 0 35 0 0 101 2
355 428
355 167
1 0 43 0 0 4096 0 36 0 0 98 2
327 429
327 351
2 0 42 0 0 4096 0 36 0 0 102 2
309 429
309 121
1 0 60 0 0 4096 0 37 0 0 97 2
282 429
282 401
2 0 25 0 0 4096 0 37 0 0 103 2
264 429
264 73
4 1 70 0 0 8320 0 41 15 0 0 5
216 532
229 532
229 1158
287 1158
287 1139
3 2 71 0 0 8320 0 38 41 0 0 5
205 473
205 500
136 500
136 541
150 541
3 1 72 0 0 4224 0 39 41 0 0 5
156 474
156 505
141 505
141 532
150 532
1 0 43 0 0 0 0 38 0 0 98 2
214 428
214 351
2 0 59 0 0 0 0 38 0 0 101 2
196 428
196 167
1 0 60 0 0 0 0 39 0 0 97 2
165 429
165 401
2 0 42 0 0 0 0 39 0 0 102 2
147 429
147 121
3 1 73 0 0 4224 0 40 16 0 0 4
106 473
106 1158
149 1158
149 1140
2 0 59 0 0 0 0 40 0 0 101 2
97 428
97 167
1 0 60 0 0 0 0 40 0 0 97 2
115 428
115 401
1 0 60 0 0 4224 0 1 0 0 0 2
72 401
1552 401
1 0 43 0 0 4224 0 2 0 0 0 2
72 351
1552 351
1 0 26 0 0 4224 0 3 0 0 0 2
72 302
1551 302
1 0 6 0 0 4224 0 4 0 0 0 2
72 254
1551 254
1 0 59 0 0 4224 0 5 0 0 0 2
69 167
1551 167
1 0 42 0 0 4224 0 6 0 0 0 2
69 121
1551 121
1 0 25 0 0 4224 0 7 0 0 0 2
69 73
1552 73
1 0 5 0 0 4224 0 8 0 0 0 2
70 32
1552 32
16
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1491 1069 1536 1084
1506 1080 1520 1091
2 S7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1361 1061 1406 1076
1376 1072 1390 1083
2 S6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1150 1062 1195 1077
1165 1074 1179 1085
2 S5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
922 1064 965 1079
936 1075 950 1086
2 S4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
665 1063 708 1078
679 1075 693 1086
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
395 1060 440 1075
410 1071 424 1082
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
262 1060 307 1075
277 1071 291 1082
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
127 1057 170 1072
141 1069 155 1080
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
10 377 47 401
20 385 36 401
2 B0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
10 332 47 356
20 340 36 356
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
12 283 49 307
22 291 38 307
2 B2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
11 230 48 254
21 238 37 254
2 B3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
8 144 45 168
18 152 34 168
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
8 99 45 123
18 107 34 123
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
7 51 44 75
17 59 33 75
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
7 10 44 34
17 18 33 34
2 A3
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
