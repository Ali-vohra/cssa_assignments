CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
17
13 Logic Switch~
5 89 468 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43355.1 0
0
13 Logic Switch~
5 90 425 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
43355.1 0
0
13 Logic Switch~
5 90 381 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
43355.1 0
0
13 Logic Switch~
5 89 335 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3421 0 0
2
43355.1 0
0
13 Logic Switch~
5 88 287 0 1 11
0 16
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8157 0 0
2
43355.1 0
0
13 Logic Switch~
5 88 239 0 1 11
0 17
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5572 0 0
2
43355.1 0
0
13 Logic Switch~
5 88 192 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8901 0 0
2
43355.1 0
0
13 Logic Switch~
5 89 145 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7361 0 0
2
43355.1 0
0
8 2-In OR~
219 643 351 0 3 22
0 5 4 2
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
4747 0 0
2
43355.1 0
0
8 2-In OR~
219 644 300 0 3 22
0 7 6 3
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
972 0 0
2
43355.1 0
0
14 Logic Display~
6 876 357 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3472 0 0
2
43355.1 0
0
14 Logic Display~
6 875 296 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9998 0 0
2
43355.1 0
0
14 Logic Display~
6 875 235 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3536 0 0
2
43355.1 0
0
9 Inverter~
13 460 505 0 2 22
0 11 10
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
4597 0 0
2
43355.1 0
0
9 2-In AND~
219 652 250 0 3 22
0 9 10 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3835 0 0
2
43355.1 0
0
8 4-2 ENC~
94 399 98 0 7 15
0 19 18 17 16 9 5 7
8 4-2 ENC~
1 0 560 0
0
2 U1
-3 -77 11 -69
0
0
0
0
0
0
15

0 3 4 5 6 9 12 13 3 4
5 6 9 12 13 0
0 0 0 0 1 0 0 0
1 U
3670 0 0
2
43355.1 0
0
8 4-2 ENC~
94 396 451 0 7 15
0 15 14 13 12 11 4 6
8 4-2 ENC~
2 0 560 0
0
2 U2
-3 -77 11 -69
0
0
0
0
0
0
15

0 3 4 5 6 9 12 13 3 4
5 6 9 12 13 0
0 0 0 0 1 0 0 0
1 U
5616 0 0
2
43355.1 0
0
18
3 1 2 0 0 4224 0 9 11 0 0 5
676 351
864 351
864 383
876 383
876 375
3 1 3 0 0 4224 0 10 12 0 0 5
677 300
863 300
863 322
875 322
875 314
6 2 4 0 0 4224 0 17 9 0 0 4
446 464
617 464
617 360
630 360
6 1 5 0 0 8320 0 16 9 0 0 4
449 111
617 111
617 342
630 342
7 2 6 0 0 4224 0 17 10 0 0 4
446 451
623 451
623 309
631 309
7 1 7 0 0 8320 0 16 10 0 0 4
449 98
623 98
623 291
631 291
3 1 8 0 0 4224 0 15 13 0 0 5
673 250
863 250
863 261
875 261
875 253
5 1 9 0 0 4224 0 16 15 0 0 4
449 152
620 152
620 241
628 241
2 2 10 0 0 8320 0 14 15 0 0 4
481 505
620 505
620 259
628 259
1 5 11 0 0 4224 0 14 17 0 0 2
445 505
446 505
1 4 12 0 0 4224 0 1 17 0 0 4
101 468
346 468
346 478
354 478
1 3 13 0 0 4224 0 2 17 0 0 4
102 425
336 425
336 464
354 464
1 2 14 0 0 4224 0 3 17 0 0 4
102 381
341 381
341 451
354 451
1 1 15 0 0 4224 0 4 17 0 0 4
101 335
346 335
346 438
354 438
1 4 16 0 0 4224 0 5 16 0 0 4
100 287
334 287
334 125
357 125
1 3 17 0 0 4224 0 6 16 0 0 4
100 239
339 239
339 111
357 111
1 2 18 0 0 4224 0 7 16 0 0 4
100 192
344 192
344 98
357 98
1 1 19 0 0 4224 0 8 16 0 0 4
101 145
349 145
349 85
357 85
11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
896 341 933 365
906 349 922 365
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
898 279 935 303
908 287 924 303
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
901 216 938 240
911 224 927 240
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
34 448 71 472
44 456 60 472
2 D0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
34 403 71 427
44 411 60 427
2 D1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
34 360 71 384
44 368 60 384
2 D2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
32 316 69 340
42 324 58 340
2 D3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
34 268 71 292
44 276 60 292
2 D4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
34 220 71 244
44 228 60 244
2 D5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
35 172 72 196
45 180 61 196
2 D6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
36 122 73 146
46 130 62 146
2 D7
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
