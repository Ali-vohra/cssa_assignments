CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
70 30 30 140 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
16
13 Logic Switch~
5 93 340 0 1 11
0 2
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
43306.4 0
0
13 Logic Switch~
5 91 282 0 1 11
0 7
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
43306.4 1
0
13 Logic Switch~
5 85 149 0 1 11
0 8
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
43306.4 2
0
13 Logic Switch~
5 83 78 0 1 11
0 13
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
43306.4 3
0
9 Inverter~
13 155 323 0 2 22
0 2 6
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U3D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 3 0
1 U
8157 0 0
2
43306.4 4
0
9 Inverter~
13 155 268 0 2 22
0 7 3
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U3C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
5572 0 0
2
43306.4 5
0
5 4071~
219 360 343 0 3 22
0 3 2 14
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U2D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 512 4 4 2 0
1 U
8901 0 0
2
43306.4 6
0
9 2-In AND~
219 368 269 0 3 22
0 5 4 15
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 4 1 0
1 U
7361 0 0
2
43306.4 7
0
5 4071~
219 232 349 0 3 22
0 3 6 4
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U2C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
4747 0 0
2
43306.4 8
0
5 4071~
219 234 273 0 3 22
0 7 2 5
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U2B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
972 0 0
2
43306.4 9
0
9 Inverter~
13 154 131 0 2 22
0 8 12
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U3B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
3472 0 0
2
43306.4 10
0
9 Inverter~
13 152 60 0 2 22
0 13 9
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
9998 0 0
2
43306.4 11
0
5 4071~
219 352 57 0 3 22
0 11 10 16
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 512 4 1 2 0
1 U
3536 0 0
2
43306.4 12
0
9 2-In AND~
219 355 128 0 3 22
0 9 8 17
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 3 1 0
1 U
4597 0 0
2
43306.4 13
0
9 2-In AND~
219 244 130 0 3 22
0 9 8 10
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3835 0 0
2
43306.4 14
0
9 2-In AND~
219 244 64 0 3 22
0 13 12 11
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3670 0 0
2
43306.4 15
0
20
1 2 2 0 0 12416 0 1 7 0 0 6
105 340
215 340
215 374
334 374
334 352
347 352
2 1 3 0 0 12416 0 6 7 0 0 6
176 268
205 268
205 369
339 369
339 334
347 334
3 2 4 0 0 4224 0 9 8 0 0 4
265 349
336 349
336 278
344 278
3 1 5 0 0 4224 0 10 8 0 0 4
267 273
336 273
336 260
344 260
2 2 6 0 0 4224 0 5 9 0 0 4
176 323
211 323
211 358
219 358
2 1 3 0 0 0 0 6 9 0 0 4
176 268
201 268
201 340
219 340
1 1 2 0 0 0 0 1 5 0 0 4
105 340
132 340
132 323
140 323
1 1 7 0 0 4096 0 2 6 0 0 4
103 282
132 282
132 268
140 268
1 2 2 0 0 0 0 1 10 0 0 4
105 340
208 340
208 282
221 282
1 1 7 0 0 4224 0 2 10 0 0 4
103 282
213 282
213 264
221 264
1 2 8 0 0 4224 0 3 14 0 0 4
97 149
318 149
318 137
331 137
2 1 9 0 0 12416 0 12 14 0 0 6
173 60
216 60
216 150
323 150
323 119
331 119
3 2 10 0 0 8320 0 15 13 0 0 4
265 130
327 130
327 66
339 66
3 1 11 0 0 4224 0 16 13 0 0 4
265 64
331 64
331 48
339 48
2 2 12 0 0 8320 0 11 16 0 0 4
175 131
202 131
202 73
220 73
2 1 9 0 0 0 0 12 15 0 0 4
173 60
207 60
207 121
220 121
1 1 13 0 0 4096 0 4 12 0 0 4
95 78
129 78
129 60
137 60
1 1 8 0 0 0 0 3 11 0 0 4
97 149
131 149
131 131
139 131
1 2 8 0 0 0 0 3 15 0 0 4
97 149
212 149
212 139
220 139
1 1 13 0 0 4224 0 4 16 0 0 4
95 78
212 78
212 55
220 55
7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
174 421 315 445
184 429 304 445
15 HALF SUBTRACTOR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
457 293 542 317
467 301 531 317
8 POS Form
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
444 76 529 100
454 84 518 100
8 SOP Form
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
382 41 483 65
392 49 472 65
10 Difference
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
372 113 441 137
382 121 430 137
6 Borrow
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
386 252 487 276
396 260 476 276
10 Difference
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
389 328 458 352
399 336 447 352
6 Borrow
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
