CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
70 0 30 110 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
26
13 Logic Switch~
5 176 412 0 1 11
0 16
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43331.5 0
0
13 Logic Switch~
5 176 212 0 10 11
0 29 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
391 0 0
2
43331.5 0
0
9 2-In AND~
219 995 347 0 3 22
0 3 4 2
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
3124 0 0
2
43331.5 0
0
9 Inverter~
13 938 305 0 2 22
0 5 4
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U8B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 6 0
1 U
3421 0 0
2
43331.5 0
0
9 Inverter~
13 938 217 0 2 22
0 6 3
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U8A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 6 0
1 U
8157 0 0
2
43331.5 0
0
5 4073~
219 862 277 0 4 22
0 9 8 7 5
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 5 0
1 U
5572 0 0
2
43331.5 0
0
9 2-In AND~
219 760 232 0 3 22
0 11 10 9
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
8901 0 0
2
43331.5 0
0
5 4030~
219 684 257 0 3 22
0 13 12 10
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U6B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 4 0
1 U
7361 0 0
2
43331.5 0
0
5 4030~
219 685 206 0 3 22
0 15 14 11
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U6A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
4747 0 0
2
43331.5 0
0
9 2-In AND~
219 822 193 0 3 22
0 7 17 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
972 0 0
2
43331.5 0
0
9 Inverter~
13 763 465 0 2 22
0 8 17
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
3472 0 0
2
43331.5 0
0
9 Inverter~
13 623 188 0 2 22
0 18 7
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
9998 0 0
2
43331.5 0
0
14 Logic Display~
6 1069 201 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3536 0 0
2
43331.5 0
0
14 Logic Display~
6 1068 278 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4597 0 0
2
43331.5 0
0
14 Logic Display~
6 1068 347 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3835 0 0
2
43331.5 0
0
8 2-In OR~
219 709 406 0 3 22
0 19 20 8
0
0 0 624 270
6 74LS32
-21 -24 21 -16
3 U5A
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3670 0 0
2
43331.5 0
0
9 2-In AND~
219 744 337 0 3 22
0 13 15 19
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U4B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
5616 0 0
2
43331.5 0
0
9 2-In AND~
219 680 338 0 3 22
0 14 15 20
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U4A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
9323 0 0
2
43331.5 0
0
8 Hex Key~
166 425 99 0 11 12
0 25 26 27 28 0 0 0 0 0
9 57
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
317 0 0
2
43331.5 0
0
6 74LS83
105 551 296 0 14 29
0 28 27 26 25 24 23 22 21 16
15 14 13 12 18
0
0 0 4848 0
5 74F83
-18 -60 17 -52
2 U3
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 0 0 0 0
1 U
3108 0 0
2
43331.5 0
0
6 74LS83
105 332 300 0 14 29
0 29 16 29 16 33 32 31 30 29
24 23 22 21 38
0
0 0 4848 0
5 74F83
-18 -60 17 -52
2 U2
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 0 0 0 0
1 U
4299 0 0
2
43331.5 0
0
9 Inverter~
13 176 368 0 2 22
0 34 30
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
9672 0 0
2
43331.5 0
0
9 Inverter~
13 176 330 0 2 22
0 35 31
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
7876 0 0
2
43331.5 0
0
9 Inverter~
13 176 292 0 2 22
0 36 32
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
6369 0 0
2
43331.5 0
0
9 Inverter~
13 175 256 0 2 22
0 37 33
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
9172 0 0
2
43331.5 0
0
8 Hex Key~
166 90 100 0 11 12
0 34 35 36 37 0 0 0 0 0
9 57
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
7100 0 0
2
43331.5 0
0
48
3 1 2 0 0 4224 0 3 15 0 0 5
1016 347
1056 347
1056 373
1068 373
1068 365
2 1 3 0 0 8320 0 5 3 0 0 4
959 217
963 217
963 338
971 338
2 2 4 0 0 8320 0 4 3 0 0 4
959 305
963 305
963 356
971 356
4 1 5 0 0 4096 0 6 4 0 0 4
883 277
915 277
915 305
923 305
3 1 6 0 0 4096 0 10 5 0 0 4
843 193
915 193
915 217
923 217
4 1 5 0 0 4224 0 6 14 0 0 5
883 277
1056 277
1056 304
1068 304
1068 296
2 3 7 0 0 4224 0 12 6 0 0 5
644 188
644 490
810 490
810 286
838 286
3 2 8 0 0 12416 0 16 6 0 0 5
712 436
712 433
830 433
830 277
838 277
3 1 9 0 0 4224 0 7 6 0 0 4
781 232
830 232
830 268
838 268
3 2 10 0 0 8320 0 8 7 0 0 4
717 257
728 257
728 241
736 241
3 1 11 0 0 8320 0 9 7 0 0 4
718 206
728 206
728 223
736 223
13 2 12 0 0 4224 0 20 8 0 0 4
583 314
653 314
653 266
668 266
12 1 13 0 0 4096 0 20 8 0 0 4
583 305
650 305
650 248
668 248
11 2 14 0 0 8192 0 20 9 0 0 4
583 296
656 296
656 215
669 215
10 1 15 0 0 8192 0 20 9 0 0 4
583 287
661 287
661 197
669 197
1 9 16 0 0 4224 0 1 20 0 0 4
188 412
511 412
511 341
519 341
3 1 6 0 0 4224 0 10 13 0 0 5
843 193
1057 193
1057 227
1069 227
1069 219
2 2 17 0 0 8320 0 11 10 0 0 4
784 465
790 465
790 202
798 202
3 1 8 0 0 128 0 16 11 0 0 3
712 436
712 465
748 465
2 1 7 0 0 128 0 12 10 0 0 4
644 188
790 188
790 184
798 184
14 1 18 0 0 8320 0 20 12 0 0 4
583 341
600 341
600 188
608 188
3 1 19 0 0 8320 0 17 16 0 0 4
742 360
742 375
721 375
721 390
3 2 20 0 0 8320 0 18 16 0 0 4
678 361
678 375
703 375
703 390
12 1 13 0 0 4224 0 20 17 0 0 3
583 305
751 305
751 315
10 2 15 0 0 4224 0 20 17 0 0 3
583 287
733 287
733 315
11 1 14 0 0 4224 0 20 18 0 0 3
583 296
687 296
687 316
10 2 15 0 0 0 0 20 18 0 0 3
583 287
669 287
669 316
13 8 21 0 0 4224 0 21 20 0 0 4
364 318
511 318
511 323
519 323
12 7 22 0 0 4224 0 21 20 0 0 4
364 309
511 309
511 314
519 314
11 6 23 0 0 4224 0 21 20 0 0 4
364 300
511 300
511 305
519 305
10 5 24 0 0 4224 0 21 20 0 0 4
364 291
511 291
511 296
519 296
1 4 25 0 0 4224 0 19 20 0 0 3
434 123
434 287
519 287
2 3 26 0 0 4224 0 19 20 0 0 3
428 123
428 278
519 278
3 2 27 0 0 4224 0 19 20 0 0 3
422 123
422 269
519 269
4 1 28 0 0 4224 0 19 20 0 0 3
416 123
416 260
519 260
1 9 29 0 0 8320 0 2 21 0 0 4
188 212
272 212
272 345
300 345
1 4 16 0 0 0 0 1 21 0 0 4
188 412
282 412
282 291
300 291
1 2 16 0 0 128 0 1 21 0 0 4
188 412
277 412
277 273
300 273
1 3 29 0 0 0 0 2 21 0 0 4
188 212
282 212
282 282
300 282
1 1 29 0 0 0 0 2 21 0 0 4
188 212
287 212
287 264
300 264
2 8 30 0 0 4224 0 22 21 0 0 4
197 368
287 368
287 327
300 327
2 7 31 0 0 4224 0 23 21 0 0 4
197 330
292 330
292 318
300 318
2 6 32 0 0 4224 0 24 21 0 0 4
197 292
287 292
287 309
300 309
2 5 33 0 0 4224 0 25 21 0 0 4
196 256
292 256
292 300
300 300
1 1 34 0 0 4224 0 26 22 0 0 3
99 124
99 368
161 368
2 1 35 0 0 4224 0 26 23 0 0 3
93 124
93 330
161 330
3 1 36 0 0 4224 0 26 24 0 0 3
87 124
87 292
161 292
4 1 37 0 0 4224 0 26 25 0 0 3
81 124
81 256
160 256
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
478 529 665 551
487 537 655 553
21 BCD COMPARATOR (10'S)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
409 37 438 59
419 45 427 61
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
75 36 102 58
84 43 92 59
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1074 338 1117 360
1083 345 1107 361
3 A>B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1075 269 1118 291
1084 276 1108 292
3 A=B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1075 188 1118 210
1084 196 1108 212
3 A<B
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
