CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
90 40 30 60 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
25
13 Logic Switch~
5 795 924 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
14 0 28 8
3 V20
10 -10 31 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5616 0 0
2
43361.9 0
0
13 Logic Switch~
5 715 923 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
14 0 28 8
3 V19
10 -10 31 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9323 0 0
2
43361.9 0
0
13 Logic Switch~
5 628 925 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
14 0 28 8
3 V18
10 -10 31 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
317 0 0
2
43361.9 0
0
13 Logic Switch~
5 540 924 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
14 0 28 8
3 V17
10 -10 31 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3108 0 0
2
43361.9 0
0
13 Logic Switch~
5 100 938 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V16
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4299 0 0
2
43361.9 0
0
13 Logic Switch~
5 101 881 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V15
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9672 0 0
2
43361.9 0
0
13 Logic Switch~
5 103 827 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V14
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7876 0 0
2
43361.9 0
0
13 Logic Switch~
5 106 776 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V13
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6369 0 0
2
43361.9 0
0
13 Logic Switch~
5 106 720 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V12
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9172 0 0
2
43361.9 0
0
13 Logic Switch~
5 108 667 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V11
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7100 0 0
2
43361.9 0
0
13 Logic Switch~
5 108 606 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V10
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3820 0 0
2
43361.9 0
0
13 Logic Switch~
5 110 547 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7678 0 0
2
43361.9 0
0
13 Logic Switch~
5 112 492 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
961 0 0
2
43361.9 0
0
13 Logic Switch~
5 113 431 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3178 0 0
2
43361.9 0
0
13 Logic Switch~
5 113 369 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3409 0 0
2
43361.9 0
0
13 Logic Switch~
5 115 306 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3951 0 0
2
43361.9 0
0
13 Logic Switch~
5 115 245 0 10 11
0 22 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8885 0 0
2
43361.9 0
0
13 Logic Switch~
5 116 185 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3780 0 0
2
43361.9 0
0
13 Logic Switch~
5 117 127 0 10 11
0 24 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9265 0 0
2
43361.9 0
0
13 Logic Switch~
5 118 72 0 10 11
0 25 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9442 0 0
2
43361.9 0
0
14 Logic Display~
6 1162 467 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9424 0 0
2
43361.9 0
0
8 2-In OR~
219 953 478 0 3 22
0 4 3 2
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
9968 0 0
2
43361.9 0
0
9 Inverter~
13 512 875 0 2 22
0 5 9
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U3A
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
9281 0 0
2
43361.9 0
0
7 74LS151
20 419 702 0 14 29
0 17 16 15 14 13 12 11 10 5
8 7 6 3 26
0
0 0 4848 0
6 74F151
-21 -60 21 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 0 0 0 0
1 U
8464 0 0
2
43361.9 0
0
7 74LS151
20 423 285 0 14 29
0 25 24 23 22 21 20 19 18 9
8 7 6 4 27
0
0 0 4848 0
6 74F151
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 0 0 0 0
1 U
7168 0 0
2
43361.9 0
0
28
3 1 2 0 0 4224 0 22 21 0 0 5
986 478
1150 478
1150 493
1162 493
1162 485
13 2 3 0 0 4224 0 24 22 0 0 4
451 729
932 729
932 487
940 487
13 1 4 0 0 4224 0 25 22 0 0 4
455 312
932 312
932 469
940 469
1 9 5 0 0 4224 0 4 24 0 0 3
541 911
541 675
457 675
1 12 6 0 0 8192 0 1 24 0 0 3
796 911
796 702
451 702
1 11 7 0 0 8192 0 2 24 0 0 3
716 910
716 693
451 693
1 10 8 0 0 4096 0 3 24 0 0 3
629 912
629 684
451 684
1 12 6 0 0 4224 0 1 25 0 0 3
796 911
796 285
455 285
1 11 7 0 0 4224 0 2 25 0 0 3
716 910
716 276
455 276
1 10 8 0 0 4224 0 3 25 0 0 3
629 912
629 267
455 267
2 9 9 0 0 4224 0 23 25 0 0 3
515 857
515 258
461 258
1 1 5 0 0 0 0 4 23 0 0 4
541 911
541 901
515 901
515 893
1 8 10 0 0 4224 0 5 24 0 0 4
112 938
364 938
364 738
387 738
1 7 11 0 0 4224 0 6 24 0 0 4
113 881
379 881
379 729
387 729
1 6 12 0 0 4224 0 7 24 0 0 4
115 827
369 827
369 720
387 720
1 5 13 0 0 4224 0 8 24 0 0 4
118 776
374 776
374 711
387 711
1 4 14 0 0 4224 0 9 24 0 0 4
118 720
379 720
379 702
387 702
1 3 15 0 0 4224 0 10 24 0 0 4
120 667
369 667
369 693
387 693
1 2 16 0 0 4224 0 11 24 0 0 4
120 606
374 606
374 684
387 684
1 1 17 0 0 4224 0 12 24 0 0 4
122 547
379 547
379 675
387 675
1 8 18 0 0 4224 0 13 25 0 0 4
124 492
373 492
373 321
391 321
1 7 19 0 0 4224 0 14 25 0 0 4
125 431
383 431
383 312
391 312
1 6 20 0 0 4224 0 15 25 0 0 4
125 369
378 369
378 303
391 303
1 5 21 0 0 4224 0 16 25 0 0 4
127 306
383 306
383 294
391 294
1 4 22 0 0 4224 0 17 25 0 0 4
127 245
368 245
368 285
391 285
1 3 23 0 0 4224 0 18 25 0 0 4
128 185
373 185
373 276
391 276
1 2 24 0 0 4224 0 19 25 0 0 4
129 127
378 127
378 267
391 267
1 1 25 0 0 4224 0 20 25 0 0 4
130 72
383 72
383 258
391 258
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
