CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
16
13 Logic Switch~
5 110 39 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3536 0 0
2
43354.9 0
0
13 Logic Switch~
5 109 114 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4597 0 0
2
43354.9 0
0
13 Logic Switch~
5 109 200 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3835 0 0
2
43354.9 1
0
13 Logic Switch~
5 109 280 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3670 0 0
2
43354.9 0
0
5 4073~
219 441 532 0 4 22
0 11 2 10 6
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 4 0
1 U
5616 0 0
2
43354.9 0
0
5 4073~
219 442 469 0 4 22
0 11 2 12 7
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 2 0
1 U
9323 0 0
2
43354.9 0
0
5 4073~
219 442 410 0 4 22
0 13 2 10 8
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 2 0
1 U
317 0 0
2
43354.9 0
0
5 4073~
219 443 353 0 4 22
0 13 2 12 9
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 2 0
1 U
3108 0 0
2
43354.9 0
0
9 2-In AND~
219 257 78 0 3 22
0 4 3 2
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
4299 0 0
2
43354.9 0
0
9 Inverter~
13 179 39 0 2 22
0 5 4
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
9672 0 0
2
43354.9 0
0
9 Inverter~
13 180 224 0 2 22
0 13 11
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
7876 0 0
2
43354.9 11
0
9 Inverter~
13 179 307 0 2 22
0 12 10
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
6369 0 0
2
43354.9 10
0
14 Logic Display~
6 818 334 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9172 0 0
2
43354.9 5
0
14 Logic Display~
6 819 391 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7100 0 0
2
43354.9 4
0
14 Logic Display~
6 818 455 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3820 0 0
2
43354.9 3
0
14 Logic Display~
6 818 516 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7678 0 0
2
43354.9 2
0
26
2 3 2 0 0 8192 0 5 9 0 0 3
417 532
278 532
278 78
2 0 2 0 0 0 0 6 0 0 5 3
418 469
312 469
312 78
2 0 2 0 0 0 0 7 0 0 5 3
418 410
345 410
345 78
2 0 2 0 0 0 0 8 0 0 5 3
419 353
380 353
380 78
3 0 2 0 0 4224 0 9 0 0 0 2
278 78
822 78
1 2 3 0 0 4224 0 2 9 0 0 3
121 114
233 114
233 87
2 1 4 0 0 4224 0 10 9 0 0 3
200 39
233 39
233 69
1 1 5 0 0 4224 0 1 10 0 0 2
122 39
164 39
4 1 6 0 0 4240 0 5 16 0 0 5
462 532
806 532
806 542
818 542
818 534
4 1 7 0 0 4240 0 6 15 0 0 5
463 469
806 469
806 481
818 481
818 473
4 1 8 0 0 4240 0 7 14 0 0 5
463 410
807 410
807 417
819 417
819 409
4 1 9 0 0 4240 0 8 13 0 0 5
464 353
806 353
806 360
818 360
818 352
3 0 10 0 0 8208 0 5 0 0 21 3
417 541
271 541
271 307
1 0 11 0 0 8208 0 5 0 0 24 3
417 523
286 523
286 224
3 0 12 0 0 8208 0 6 0 0 23 3
418 478
303 478
303 280
1 0 11 0 0 16 0 6 0 0 24 3
418 460
320 460
320 224
3 0 10 0 0 16 0 7 0 0 21 3
418 419
337 419
337 307
1 0 13 0 0 8208 0 7 0 0 26 3
418 401
354 401
354 200
3 0 12 0 0 16 0 8 0 0 23 3
419 362
371 362
371 280
1 0 13 0 0 16 0 8 0 0 26 3
419 344
390 344
390 200
2 0 10 0 0 4240 0 12 0 0 0 2
200 307
824 307
1 1 12 0 0 16 0 4 12 0 0 4
121 280
156 280
156 307
164 307
1 0 12 0 0 4240 0 4 0 0 0 2
121 280
822 280
2 0 11 0 0 4240 0 11 0 0 0 2
201 224
822 224
1 1 13 0 0 16 0 3 11 0 0 4
121 200
157 200
157 224
165 224
1 0 13 0 0 4240 0 3 0 0 0 2
121 200
822 200
8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
51 90 88 114
61 98 77 114
2 E1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
49 18 86 42
59 26 75 42
2 E2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
849 499 886 523
859 507 875 523
2 D0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
850 440 887 464
860 448 876 464
2 D1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
849 375 886 399
859 383 875 399
2 D2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
850 318 887 342
860 326 876 342
2 D3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
54 259 91 283
64 267 80 283
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
53 176 90 200
63 184 79 200
2 A1
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
