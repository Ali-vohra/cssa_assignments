CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
110 60 30 110 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
15
13 Logic Switch~
5 144 470 0 1 11
0 7
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 142 388 0 1 11
0 6
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 127 216 0 1 11
0 8
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 128 150 0 1 11
0 9
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 391 412 0 3 22
0 2 3 14
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 4 1 0
1 U
8157 0 0
2
5.89855e-315 0
0
9 Inverter~
13 203 457 0 2 22
0 7 4
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
5572 0 0
2
5.89855e-315 0
0
9 Inverter~
13 202 402 0 2 22
0 6 5
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
8901 0 0
2
5.89855e-315 0
0
5 4071~
219 273 456 0 3 22
0 5 4 3
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 3 0
1 U
7361 0 0
2
5.89855e-315 0
0
5 4071~
219 268 387 0 3 22
0 6 7 2
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 3 0
1 U
4747 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 330 287 0 3 22
0 9 8 15
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 3 1 0
1 U
972 0 0
2
5.89855e-315 0
0
5 4071~
219 416 167 0 3 22
0 11 10 16
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 512 4 1 3 0
1 U
3472 0 0
2
5.89855e-315 0
0
9 Inverter~
13 257 166 0 2 22
0 9 12
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
9998 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 330 209 0 3 22
0 8 12 10
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3536 0 0
2
5.89855e-315 0
0
9 Inverter~
13 258 213 0 2 22
0 8 13
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
4597 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 332 141 0 3 22
0 9 13 11
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3835 0 0
2
5.89855e-315 0
0
19
3 0 2 0 0 4224 0 9 0 0 0 3
301 387
301 514
413 514
3 2 3 0 0 4224 0 8 5 0 0 4
306 456
359 456
359 421
367 421
3 1 2 0 0 0 0 9 5 0 0 4
301 387
359 387
359 403
367 403
2 2 4 0 0 4224 0 6 8 0 0 4
224 457
252 457
252 465
260 465
2 1 5 0 0 8320 0 7 8 0 0 4
223 402
250 402
250 447
260 447
1 1 6 0 0 4096 0 2 7 0 0 4
154 388
179 388
179 402
187 402
1 1 7 0 0 4096 0 1 6 0 0 4
156 470
180 470
180 457
188 457
1 2 7 0 0 4224 0 1 9 0 0 4
156 470
247 470
247 396
255 396
1 1 6 0 0 4224 0 2 9 0 0 4
154 388
247 388
247 378
255 378
1 2 8 0 0 4096 0 3 10 0 0 4
139 216
229 216
229 296
306 296
1 1 9 0 0 4096 0 4 10 0 0 4
140 150
288 150
288 278
306 278
3 2 10 0 0 4224 0 13 11 0 0 4
351 209
395 209
395 176
403 176
3 1 11 0 0 4224 0 15 11 0 0 4
353 141
395 141
395 158
403 158
2 2 12 0 0 8320 0 12 13 0 0 4
278 166
298 166
298 218
306 218
1 1 9 0 0 0 0 4 12 0 0 4
140 150
234 150
234 166
242 166
1 1 8 0 0 4224 0 3 13 0 0 4
139 216
239 216
239 200
306 200
2 2 13 0 0 8320 0 14 15 0 0 4
279 213
295 213
295 150
308 150
1 1 8 0 0 0 0 3 14 0 0 4
139 216
235 216
235 213
243 213
1 1 9 0 0 4224 0 4 15 0 0 4
140 150
300 150
300 132
308 132
7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
231 553 326 577
238 559 318 575
10 HALF ADDER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
451 149 496 173
461 157 485 173
3 Sum
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
348 271 409 295
358 279 398 295
5 Carry
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
233 67 318 91
243 75 307 91
8 SOP Form
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
410 396 455 420
420 404 444 420
3 Sum
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
409 497 470 521
419 505 459 521
5 Carry
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
225 325 310 349
235 333 299 349
8 POS Form
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
