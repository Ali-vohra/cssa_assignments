CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
14
13 Logic Switch~
5 71 94 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43335 0
0
13 Logic Switch~
5 69 228 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
43335 0
0
13 Logic Switch~
5 70 177 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
43335 0
0
13 Logic Switch~
5 72 51 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3421 0 0
2
43335 0
0
14 Logic Display~
6 504 443 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8157 0 0
2
43335.1 0
0
14 Logic Display~
6 416 445 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5572 0 0
2
43335.1 0
0
14 Logic Display~
6 301 447 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8901 0 0
2
43335.1 0
0
14 Logic Display~
6 159 450 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7361 0 0
2
43335.1 0
0
9 2-In AND~
219 350 278 0 3 22
0 2 3 10
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1D
-13 -12 8 -4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
4747 0 0
2
43335.1 0
0
9 2-In AND~
219 242 277 0 3 22
0 2 4 11
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1C
-12 -11 9 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
972 0 0
2
43335.1 0
0
9 2-In AND~
219 202 277 0 3 22
0 5 3 12
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1B
-12 -11 9 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3472 0 0
2
43335.1 0
0
9 2-In AND~
219 133 276 0 3 22
0 5 4 13
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1A
-12 -11 9 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
9998 0 0
2
43335.1 0
0
2 HA
94 220 354 0 4 9
0 11 12 8 9
2 HA
1 0 656 0
0
2 U2
-7 -28 7 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 U
3536 0 0
2
43334.7 0
0
2 HA
94 346 353 0 4 9
0 8 10 6 7
2 HA
2 0 656 0
0
2 U3
-7 -28 7 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 U
4597 0 0
2
43334.7 0
0
20
1 0 2 0 0 4096 0 9 0 0 10 2
357 256
357 177
2 0 3 0 0 4096 0 9 0 0 12 2
339 256
339 51
1 0 2 0 0 0 0 10 0 0 10 2
249 255
249 177
2 0 4 0 0 4096 0 10 0 0 11 2
231 255
231 94
1 0 5 0 0 4096 0 11 0 0 9 2
209 255
209 228
2 0 3 0 0 0 0 11 0 0 12 2
191 255
191 51
1 0 5 0 0 0 0 12 0 0 9 2
140 254
140 228
2 0 4 0 0 0 0 12 0 0 11 2
122 254
122 94
1 0 5 0 0 4224 0 2 0 0 0 2
81 228
523 228
1 0 2 0 0 4224 0 3 0 0 0 2
82 177
523 177
1 0 4 0 0 4224 0 1 0 0 0 2
83 94
524 94
1 0 3 0 0 4224 0 4 0 0 0 2
84 51
524 51
3 1 6 0 0 8320 0 14 5 0 0 5
379 362
472 362
472 479
504 479
504 461
4 1 7 0 0 8320 0 14 6 0 0 5
379 353
394 353
394 478
416 478
416 463
3 1 8 0 0 4224 0 13 14 0 0 4
253 363
283 363
283 353
313 353
4 1 9 0 0 8320 0 13 7 0 0 5
253 354
274 354
274 477
301 477
301 465
3 2 10 0 0 8320 0 9 14 0 0 4
348 301
291 301
291 362
313 362
3 1 11 0 0 8320 0 10 13 0 0 5
240 300
240 311
169 311
169 354
187 354
3 2 12 0 0 8320 0 11 13 0 0 4
200 300
160 300
160 363
187 363
3 1 13 0 0 4224 0 12 8 0 0 4
131 299
131 477
159 477
159 468
8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
490 501 527 525
500 509 516 525
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
398 501 435 525
408 509 424 525
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
284 500 321 524
294 508 310 524
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
141 501 178 525
151 509 167 525
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
14 204 51 228
24 212 40 228
2 B0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
15 156 52 180
25 164 41 180
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
16 75 53 99
26 83 42 99
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
18 32 55 56
28 40 44 56
2 A1
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
