CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
180 70 30 110 10
176 80 1534 843
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
24
13 Logic Switch~
5 536 191 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89857e-315 0
0
13 Logic Switch~
5 332 301 0 1 11
0 22
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
43319.7 0
0
5 4049~
219 645 679 0 2 22
0 4 3
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 1 0
1 U
3124 0 0
2
43319.7 0
0
5 4081~
219 716 709 0 3 22
0 3 5 2
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U8A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
3421 0 0
2
43319.7 0
0
9 2-In AND~
219 634 634 0 3 22
0 5 6 4
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
8157 0 0
2
43319.7 0
0
5 4082~
219 548 565 0 5 22
0 10 9 8 7 6
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U6A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 4 0
1 U
5572 0 0
2
43319.7 0
0
14 Logic Display~
6 986 711 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8901 0 0
2
43319.7 0
0
14 Logic Display~
6 983 623 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7361 0 0
2
43319.7 0
0
14 Logic Display~
6 980 539 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4747 0 0
2
43319.7 0
0
9 Inverter~
13 462 362 0 2 22
0 11 5
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
972 0 0
2
5.89857e-315 0
0
5 4030~
219 536 497 0 3 22
0 7 5 13
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U4D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 2 0
1 U
3472 0 0
2
5.89857e-315 0
0
5 4030~
219 539 445 0 3 22
0 8 5 14
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U4C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
9998 0 0
2
5.89857e-315 5.26354e-315
0
5 4030~
219 541 394 0 3 22
0 9 5 15
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U4B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
3536 0 0
2
5.89857e-315 0
0
5 4030~
219 539 341 0 3 22
0 10 5 16
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U4A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
4597 0 0
2
5.89857e-315 0
0
14 Logic Display~
6 968 297 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3835 0 0
2
43319.7 1
0
12 Hex Display~
7 861 160 0 18 19
10 18 19 20 21 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3670 0 0
2
43319.7 2
0
6 74LS83
105 643 270 0 14 29
0 16 15 14 13 12 12 12 12 11
21 20 19 18 17
0
0 0 4848 0
7 74LS83A
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
5616 0 0
2
43319.7 3
0
5 4049~
219 265 449 0 2 22
0 24 23
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 1 0
1 U
9323 0 0
2
43319.7 4
0
5 4049~
219 265 410 0 2 22
0 26 25
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 1 0
1 U
317 0 0
2
43319.7 5
0
5 4049~
219 267 371 0 2 22
0 28 27
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 1 0
1 U
3108 0 0
2
43319.7 6
0
5 4049~
219 267 333 0 2 22
0 30 29
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 1 0
1 U
4299 0 0
2
43319.7 7
0
8 Hex Key~
166 205 170 0 11 12
0 24 26 28 30 0 0 0 0 0
6 54
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
9672 0 0
2
43319.7 8
0
8 Hex Key~
166 310 171 0 11 12
0 31 32 33 34 0 0 0 0 0
5 53
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
7876 0 0
2
43319.7 9
0
6 74LS83
105 451 273 0 14 29
0 34 33 32 31 29 27 25 23 22
10 9 8 7 11
0
0 0 4848 0
7 74LS83A
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
6369 0 0
2
43319.7 10
0
48
3 1 2 0 0 4224 0 4 7 0 0 5
737 709
974 709
974 737
986 737
986 729
2 1 3 0 0 8320 0 3 4 0 0 4
666 679
679 679
679 700
692 700
3 1 4 0 0 8192 0 5 3 0 0 6
655 634
670 634
670 694
622 694
622 679
630 679
2 2 5 0 0 8320 0 10 4 0 0 4
483 362
684 362
684 718
692 718
3 1 4 0 0 4224 0 5 8 0 0 5
655 634
971 634
971 649
983 649
983 641
5 2 6 0 0 8320 0 6 5 0 0 4
569 565
597 565
597 643
610 643
2 1 5 0 0 128 0 10 5 0 0 4
483 362
602 362
602 625
610 625
4 13 7 0 0 8320 0 6 24 0 0 4
524 579
516 579
516 291
483 291
12 3 8 0 0 8320 0 24 6 0 0 4
483 282
491 282
491 570
524 570
2 11 9 0 0 8320 0 6 24 0 0 4
524 561
516 561
516 273
483 273
10 1 10 0 0 8320 0 24 6 0 0 4
483 264
491 264
491 552
524 552
14 1 11 0 0 12416 0 24 9 0 0 5
483 318
607 318
607 565
980 565
980 557
8 1 12 0 0 8320 0 17 1 0 0 4
611 297
562 297
562 191
548 191
1 7 12 0 0 0 0 1 17 0 0 4
548 191
593 191
593 288
611 288
6 1 12 0 0 0 0 17 1 0 0 4
611 279
557 279
557 191
548 191
1 5 12 0 0 0 0 1 17 0 0 4
548 191
598 191
598 270
611 270
14 9 11 0 0 128 0 24 17 0 0 4
483 318
598 318
598 315
611 315
4 3 13 0 0 8320 0 17 11 0 0 4
611 261
579 261
579 497
569 497
3 3 14 0 0 8320 0 17 12 0 0 4
611 252
585 252
585 445
572 445
2 3 15 0 0 8320 0 17 13 0 0 4
611 243
582 243
582 394
574 394
3 1 16 0 0 8320 0 14 17 0 0 4
572 341
603 341
603 234
611 234
2 2 5 0 0 128 0 10 11 0 0 4
483 362
487 362
487 506
520 506
2 2 5 0 0 0 0 10 12 0 0 4
483 362
490 362
490 454
523 454
2 2 5 0 0 0 0 10 13 0 0 4
483 362
497 362
497 403
525 403
2 2 5 0 0 0 0 10 14 0 0 4
483 362
515 362
515 350
523 350
14 1 11 0 0 0 0 24 10 0 0 6
483 318
487 318
487 377
439 377
439 362
447 362
13 1 7 0 0 128 0 24 11 0 0 4
483 291
502 291
502 488
520 488
12 1 8 0 0 128 0 24 12 0 0 4
483 282
505 282
505 436
523 436
11 1 9 0 0 128 0 24 13 0 0 4
483 273
512 273
512 385
525 385
10 1 10 0 0 128 0 24 14 0 0 4
483 264
515 264
515 332
523 332
14 1 17 0 0 4224 0 17 15 0 0 5
675 315
956 315
956 323
968 323
968 315
13 1 18 0 0 4224 0 17 16 0 0 3
675 288
870 288
870 184
12 2 19 0 0 4224 0 17 16 0 0 3
675 279
864 279
864 184
11 3 20 0 0 4224 0 17 16 0 0 3
675 270
858 270
858 184
10 4 21 0 0 4224 0 17 16 0 0 3
675 261
852 261
852 184
1 9 22 0 0 4224 0 2 24 0 0 4
344 301
391 301
391 318
419 318
2 8 23 0 0 8320 0 18 24 0 0 4
286 449
396 449
396 300
419 300
1 1 24 0 0 4224 0 22 18 0 0 3
214 194
214 449
250 449
2 7 25 0 0 8320 0 19 24 0 0 4
286 410
401 410
401 291
419 291
2 1 26 0 0 4224 0 22 19 0 0 3
208 194
208 410
250 410
2 6 27 0 0 4224 0 20 24 0 0 4
288 371
406 371
406 282
419 282
3 1 28 0 0 4224 0 22 20 0 0 3
202 194
202 371
252 371
2 5 29 0 0 4224 0 21 24 0 0 4
288 333
411 333
411 273
419 273
4 1 30 0 0 4224 0 22 21 0 0 3
196 194
196 333
252 333
1 4 31 0 0 8320 0 23 24 0 0 3
319 195
319 264
419 264
2 3 32 0 0 8320 0 23 24 0 0 3
313 195
313 255
419 255
3 2 33 0 0 8320 0 23 24 0 0 3
307 195
307 246
419 246
4 1 34 0 0 8320 0 23 24 0 0 3
301 195
301 237
419 237
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
501 99 696 121
510 106 686 122
22 4 BIT COMPARATOR (1'S)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
996 702 1039 724
1005 709 1029 725
3 A<B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
995 610 1038 632
1004 617 1028 633
3 A=B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
994 532 1031 556
1000 537 1024 553
3 A>B
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
