CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 90 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
22
13 Logic Switch~
5 278 83 0 1 11
0 2
0
0 0 21344 270
2 0V
-6 -21 8 -13
2 V5
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 168 86 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 126 86 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3124 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 83 86 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 45 86 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8157 0 0
2
5.89859e-315 0
0
14 Logic Display~
6 1172 580 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5572 0 0
2
5.89859e-315 0
0
14 Logic Display~
6 1170 506 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8901 0 0
2
5.89859e-315 0
0
6 74LS83
105 801 376 0 14 29
0 2 2 4 7 2 2 2 6 2
24 25 3 5 26
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U5
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
7361 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 207 430 0 3 22
0 6 10 9
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U4B
-13 -2 8 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
4747 0 0
2
5.89859e-315 0
0
14 Logic Display~
6 1169 432 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
972 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 207 381 0 3 22
0 6 14 13
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U4A
-13 -4 8 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3472 0 0
2
5.89859e-315 0
0
14 Logic Display~
6 1168 363 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9998 0 0
2
5.89859e-315 0
0
6 74LS83
105 633 288 0 14 29
0 2 9 12 16 2 8 2 10 2
4 7 11 15 27
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U3
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
3536 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 208 311 0 3 22
0 10 14 18
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U1D
-13 -4 8 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
4597 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 208 260 0 3 22
0 6 20 19
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U1C
-13 -3 8 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3835 0 0
2
5.89859e-315 0
0
14 Logic Display~
6 1167 290 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3670 0 0
2
5.89859e-315 0
0
14 Logic Display~
6 1165 218 0 1 2
10 21
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5616 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 209 203 0 3 22
0 10 20 22
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U1B
-13 -4 8 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
9323 0 0
2
5.89859e-315 0
0
6 74LS83
105 438 201 0 14 29
0 13 19 22 23 2 18 2 14 2
12 16 17 21 8
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U2
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
317 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 209 159 0 3 22
0 14 20 23
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U1A
-13 -4 8 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3108 0 0
2
5.89859e-315 0
0
14 Logic Display~
6 1164 157 0 1 2
10 28
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 1 0 0 0
1 L
4299 0 0
2
5.89859e-315 0
0
14 Logic Display~
6 1162 97 0 1 2
10 20
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9672 0 0
2
5.89859e-315 0
0
50
0 1 2 0 0 8192 0 0 8 2 0 3
724 349
724 340
769 340
0 2 2 0 0 8192 0 0 8 3 0 3
714 376
714 349
769 349
0 5 2 0 0 8192 0 0 8 4 0 3
704 385
704 376
769 376
0 6 2 0 0 8192 0 0 8 11 0 3
691 421
691 385
769 385
12 1 3 0 0 4224 0 8 6 0 0 5
833 385
1110 385
1110 608
1172 608
1172 598
0 7 2 0 0 0 0 0 8 11 0 3
735 421
735 394
769 394
10 3 4 0 0 4224 0 13 8 0 0 4
665 279
756 279
756 358
769 358
0 1 2 0 0 0 0 0 13 9 0 3
562 288
562 252
601 252
0 5 2 0 0 0 0 0 13 20 0 3
546 306
546 288
601 288
13 1 5 0 0 4224 0 8 7 0 0 5
833 394
1120 394
1120 534
1170 534
1170 524
0 9 2 0 0 8192 0 0 8 18 0 3
554 333
554 421
769 421
8 0 6 0 0 12416 0 8 0 0 50 4
769 403
664 403
664 473
45 473
11 4 7 0 0 4224 0 13 8 0 0 4
665 288
761 288
761 367
769 367
14 6 8 0 0 4224 0 19 13 0 0 4
470 246
578 246
578 297
601 297
3 2 9 0 0 4224 0 9 13 0 0 4
228 430
583 430
583 261
601 261
2 0 10 0 0 4096 0 9 0 0 49 2
183 439
83 439
1 0 6 0 0 0 0 9 0 0 50 2
183 421
45 421
0 9 2 0 0 0 0 0 13 20 0 3
513 306
513 333
601 333
12 1 11 0 0 4224 0 13 10 0 0 5
665 297
1131 297
1131 459
1169 459
1169 450
0 7 2 0 0 8320 0 0 13 41 0 3
330 246
330 306
601 306
10 3 12 0 0 4224 0 19 13 0 0 4
470 192
588 192
588 270
601 270
1 5 2 0 0 0 0 1 19 0 0 3
278 95
278 201
406 201
3 1 13 0 0 8320 0 11 19 0 0 4
228 381
380 381
380 165
406 165
2 0 14 0 0 4096 0 11 0 0 48 2
183 390
126 390
1 0 6 0 0 0 0 11 0 0 50 2
183 372
45 372
13 1 15 0 0 4224 0 13 12 0 0 4
665 306
1140 306
1140 381
1168 381
8 0 10 0 0 12288 0 13 0 0 49 4
601 315
405 315
405 351
83 351
11 4 16 0 0 4224 0 19 13 0 0 4
470 201
593 201
593 279
601 279
12 1 17 0 0 4224 0 19 16 0 0 5
470 210
1148 210
1148 316
1167 316
1167 308
3 6 18 0 0 4224 0 14 19 0 0 4
229 311
398 311
398 210
406 210
3 2 19 0 0 4224 0 15 19 0 0 4
229 260
388 260
388 174
406 174
2 0 14 0 0 4096 0 14 0 0 48 2
184 320
126 320
1 0 10 0 0 0 0 14 0 0 49 2
184 302
83 302
2 0 20 0 0 4096 0 15 0 0 47 2
184 269
168 269
1 0 6 0 0 0 0 15 0 0 50 2
184 251
45 251
13 1 21 0 0 4224 0 19 17 0 0 5
470 219
1153 219
1153 244
1165 244
1165 236
1 7 2 0 0 0 0 1 19 0 0 3
278 95
278 219
406 219
3 3 22 0 0 4224 0 18 19 0 0 4
230 203
392 203
392 183
406 183
2 0 20 0 0 4096 0 18 0 0 47 2
185 212
168 212
1 0 10 0 0 0 0 18 0 0 49 2
185 194
83 194
1 9 2 0 0 0 0 1 19 0 0 3
278 95
278 246
406 246
8 0 14 0 0 4096 0 19 0 0 48 2
406 228
126 228
3 4 23 0 0 4224 0 20 19 0 0 4
230 159
398 159
398 192
406 192
2 0 20 0 0 0 0 20 0 0 47 2
185 168
168 168
1 0 14 0 0 0 0 20 0 0 48 2
185 150
126 150
0 1 20 0 0 4224 0 0 22 47 0 3
168 114
1162 114
1162 115
1 0 20 0 0 0 0 2 0 0 0 2
168 98
168 601
1 0 14 0 0 4224 0 3 0 0 0 2
126 98
126 600
1 0 10 0 0 4224 0 4 0 0 0 2
83 98
83 601
1 0 6 0 0 0 0 5 0 0 0 2
45 98
45 600
12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
28 14 65 38
38 22 54 38
2 A3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
66 14 103 38
76 22 92 38
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
108 15 145 39
118 23 134 39
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
151 15 188 39
161 23 177 39
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1174 82 1211 106
1184 90 1200 106
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1175 143 1212 167
1185 151 1201 167
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1175 203 1212 227
1185 211 1201 227
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1176 275 1213 299
1186 283 1202 299
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1177 346 1214 370
1187 354 1203 370
2 S4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1177 415 1214 439
1187 423 1203 439
2 S5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1177 491 1214 515
1187 499 1203 515
2 S6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1179 566 1216 590
1189 574 1205 590
2 S7
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
