CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 279 267 0 1 11
0 10
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 576 265 0 1 11
0 11
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89855e-315 0
0
12 Hex Display~
7 664 84 0 18 19
10 2 3 4 5 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3124 0 0
2
5.89855e-315 0
0
12 Hex Display~
7 375 93 0 18 19
10 6 7 8 9 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3421 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 523 201 0 3 22
0 14 13 12
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U3C
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
8157 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 363 200 0 3 22
0 8 8 13
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U3B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
5572 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 653 200 0 3 22
0 4 3 14
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U3A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
8901 0 0
2
5.89855e-315 0
0
7 Pulser~
4 561 362 0 10 12
0 16 17 15 18 0 0 5 5 3
8
0
0 0 4640 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7361 0 0
2
5.89855e-315 0
0
6 74LS90
107 652 292 0 10 21
0 11 11 12 12 15 2 5 4 3
2
0
0 0 4832 0
6 74LS90
-21 -51 21 -43
2 U2
-7 -52 7 -44
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
4747 0 0
2
5.89855e-315 0
0
6 74LS90
107 362 295 0 10 21
0 10 10 12 12 5 6 9 8 7
6
0
0 0 4832 0
6 74LS90
-21 -51 21 -43
2 U1
-7 -52 7 -44
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
972 0 0
2
5.89855e-315 0
0
26
10 1 2 0 0 8320 0 9 3 0 0 5
684 319
718 319
718 131
673 131
673 108
9 2 3 0 0 8320 0 9 3 0 0 5
684 301
713 301
713 126
667 126
667 108
8 3 4 0 0 8320 0 9 3 0 0 5
684 283
708 283
708 121
661 121
661 108
7 4 5 0 0 8192 0 9 3 0 0 5
684 265
703 265
703 116
655 116
655 108
10 1 6 0 0 8320 0 10 4 0 0 5
394 322
433 322
433 140
384 140
384 117
9 2 7 0 0 8320 0 10 4 0 0 5
394 304
428 304
428 135
378 135
378 117
8 3 8 0 0 8320 0 10 4 0 0 5
394 286
423 286
423 130
372 130
372 117
7 4 9 0 0 8320 0 10 4 0 0 5
394 268
418 268
418 125
366 125
366 117
1 2 10 0 0 12416 0 1 10 0 0 4
291 267
306 267
306 277
330 277
1 1 10 0 0 0 0 1 10 0 0 4
291 267
311 267
311 268
330 268
1 2 11 0 0 4096 0 2 9 0 0 4
588 265
606 265
606 274
620 274
1 1 11 0 0 4224 0 2 9 0 0 2
588 265
620 265
3 4 12 0 0 12288 0 5 9 0 0 4
496 201
489 201
489 292
620 292
3 3 12 0 0 0 0 5 9 0 0 4
496 201
494 201
494 283
620 283
3 4 12 0 0 8320 0 5 10 0 0 6
496 201
413 201
413 347
306 347
306 295
330 295
3 3 12 0 0 0 0 5 10 0 0 6
496 201
408 201
408 248
316 248
316 286
330 286
3 2 13 0 0 12416 0 6 5 0 0 6
336 200
334 200
334 180
551 180
551 192
541 192
3 1 14 0 0 4224 0 7 5 0 0 4
626 200
551 200
551 210
541 210
8 2 8 0 0 0 0 10 6 0 0 4
394 286
403 286
403 191
381 191
8 1 8 0 0 0 0 10 6 0 0 4
394 286
398 286
398 209
381 209
9 2 3 0 0 0 0 9 7 0 0 4
684 301
698 301
698 191
671 191
8 1 4 0 0 0 0 9 7 0 0 4
684 283
688 283
688 209
671 209
10 6 6 0 0 0 0 10 10 0 0 6
394 322
398 322
398 342
311 342
311 322
324 322
7 5 5 0 0 12416 0 9 10 0 0 6
684 265
693 265
693 337
316 337
316 313
324 313
10 6 2 0 0 0 0 9 9 0 0 6
684 319
688 319
688 334
601 334
601 319
614 319
3 5 15 0 0 8320 0 8 9 0 0 4
585 353
606 353
606 310
614 310
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
408 401 589 425
418 409 578 425
20 DIVIDE BY 45 COUNTER
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
