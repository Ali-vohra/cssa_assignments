CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
270 290 30 160 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
12
13 Logic Switch~
5 784 163 0 1 11
0 6
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 379 291 0 1 11
0 5
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89855e-315 0
0
5 4071~
219 820 327 0 3 22
0 4 3 2
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U5A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
3124 0 0
2
5.89855e-315 0
0
12 Hex Display~
7 850 106 0 18 19
10 2 6 6 6 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3421 0 0
2
5.89855e-315 0
0
12 Hex Display~
7 911 107 0 18 19
10 7 8 9 10 0 0 0 0 0
0 1 1 1 1 1 1 1 8
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
8157 0 0
2
5.89855e-315 0
0
8 3-In OR~
219 609 399 0 4 22
0 12 3 13 11
0
0 0 608 270
4 4075
-14 -24 14 -16
3 U4A
28 -7 49 1
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 2 0
1 U
5572 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 644 342 0 3 22
0 14 15 12
0
0 0 608 270
6 74LS08
-21 -24 21 -16
3 U3B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
8901 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 574 344 0 3 22
0 16 15 13
0
0 0 608 270
6 74LS08
-21 -24 21 -16
3 U3A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
7361 0 0
2
5.89855e-315 0
0
6 74LS83
105 729 240 0 14 29
0 15 16 14 17 5 11 11 5 5
10 9 8 7 4
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U2
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
4747 0 0
2
5.89855e-315 0
0
8 Hex Key~
166 293 110 0 11 12
0 22 23 24 25 0 0 0 0 0
9 57
0
0 0 4640 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
972 0 0
2
5.89855e-315 0
0
8 Hex Key~
166 388 111 0 11 12
0 18 19 20 21 0 0 0 0 0
9 57
0
0 0 4640 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3472 0 0
2
5.89855e-315 0
0
6 74LS83
105 497 243 0 14 29
0 25 24 23 22 21 20 19 18 5
15 16 14 17 3
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
9998 0 0
2
5.89855e-315 0
0
35
3 1 2 0 0 8320 0 3 4 0 0 3
853 327
859 327
859 130
14 2 3 0 0 4224 0 12 3 0 0 4
529 288
693 288
693 336
807 336
14 1 4 0 0 4224 0 9 3 0 0 4
761 285
799 285
799 318
807 318
1 9 5 0 0 12416 0 2 9 0 0 6
391 291
446 291
446 308
674 308
674 285
697 285
1 2 6 0 0 4224 0 1 4 0 0 3
796 163
853 163
853 130
1 3 6 0 0 0 0 1 4 0 0 3
796 163
847 163
847 130
1 4 6 0 0 0 0 1 4 0 0 3
796 163
841 163
841 130
13 1 7 0 0 4224 0 9 5 0 0 3
761 258
920 258
920 131
12 2 8 0 0 4224 0 9 5 0 0 3
761 249
914 249
914 131
11 3 9 0 0 4224 0 9 5 0 0 3
761 240
908 240
908 131
10 4 10 0 0 4224 0 9 5 0 0 3
761 231
902 231
902 131
1 8 5 0 0 0 0 2 9 0 0 6
391 291
451 291
451 303
679 303
679 267
697 267
1 5 5 0 0 0 0 2 9 0 0 6
391 291
461 291
461 187
669 187
669 240
697 240
4 7 11 0 0 12288 0 6 9 0 0 5
612 429
612 431
684 431
684 258
697 258
4 6 11 0 0 12416 0 6 9 0 0 5
612 429
612 426
689 426
689 249
697 249
14 2 3 0 0 0 0 12 6 0 0 3
529 288
612 288
612 384
3 1 12 0 0 8320 0 7 6 0 0 4
642 365
642 370
621 370
621 383
3 3 13 0 0 8320 0 8 6 0 0 4
572 367
572 371
603 371
603 383
12 1 14 0 0 4096 0 12 7 0 0 3
529 252
651 252
651 320
10 2 15 0 0 4096 0 12 7 0 0 3
529 234
633 234
633 320
11 1 16 0 0 8192 0 12 8 0 0 3
529 243
581 243
581 322
10 2 15 0 0 0 0 12 8 0 0 3
529 234
563 234
563 322
13 4 17 0 0 4224 0 12 9 0 0 4
529 261
674 261
674 231
697 231
12 3 14 0 0 4224 0 12 9 0 0 4
529 252
679 252
679 222
697 222
11 2 16 0 0 4224 0 12 9 0 0 4
529 243
684 243
684 213
697 213
10 1 15 0 0 4224 0 12 9 0 0 4
529 234
689 234
689 204
697 204
1 9 5 0 0 0 0 2 12 0 0 4
391 291
457 291
457 288
465 288
1 8 18 0 0 4224 0 11 12 0 0 3
397 135
397 270
465 270
2 7 19 0 0 4224 0 11 12 0 0 3
391 135
391 261
465 261
3 6 20 0 0 4224 0 11 12 0 0 3
385 135
385 252
465 252
4 5 21 0 0 4224 0 11 12 0 0 3
379 135
379 243
465 243
1 4 22 0 0 8320 0 10 12 0 0 3
302 134
302 234
465 234
2 3 23 0 0 8320 0 10 12 0 0 3
296 134
296 225
465 225
3 2 24 0 0 8320 0 10 12 0 0 3
290 134
290 216
465 216
4 1 25 0 0 8320 0 10 12 0 0 3
284 134
284 207
465 207
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
576 462 661 486
582 467 654 483
9 BCD ADDER
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
