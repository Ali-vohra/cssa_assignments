CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
50 10 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
21
13 Logic Switch~
5 490 324 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43331.8 0
0
13 Logic Switch~
5 172 390 0 1 11
0 26
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
43331.8 0
0
13 Logic Switch~
5 173 228 0 10 11
0 27 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3124 0 0
2
43331.8 0
0
9 2-In AND~
219 857 195 0 3 22
0 4 3 2
0
0 0 624 90
6 74LS08
-21 -24 21 -16
3 U6B
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3421 0 0
2
43331.8 0
0
9 Inverter~
13 857 352 0 2 22
0 5 3
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U7A
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
8157 0 0
2
43331.8 0
0
9 Inverter~
13 854 295 0 2 22
0 6 4
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U3F
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
5572 0 0
2
43331.8 0
0
9 2-In AND~
219 795 312 0 3 22
0 8 7 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
8901 0 0
2
43331.8 0
0
5 4082~
219 658 328 0 5 22
0 12 11 10 9 8
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U5A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 2 0
1 U
7361 0 0
2
43331.8 0
0
9 Inverter~
13 682 407 0 2 22
0 5 7
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
4747 0 0
2
43331.8 0
0
14 Logic Display~
6 960 202 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
972 0 0
2
43331.8 0
0
14 Logic Display~
6 962 324 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3472 0 0
2
43331.8 0
0
14 Logic Display~
6 965 432 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9998 0 0
2
43331.8 0
0
6 74LS83
105 603 324 0 14 29
0 17 16 15 14 21 20 19 18 13
12 11 10 9 5
0
0 0 4848 0
5 74F83
-18 -60 17 -52
2 U4
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 0 0 0 0
1 U
3536 0 0
2
43331.8 0
0
9 Inverter~
13 417 478 0 2 22
0 22 18
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
4597 0 0
2
43331.8 0
0
9 Inverter~
13 416 440 0 2 22
0 23 19
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3835 0 0
2
43331.8 0
0
9 Inverter~
13 415 402 0 2 22
0 24 20
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
3670 0 0
2
43331.8 0
0
9 Inverter~
13 414 365 0 2 22
0 25 21
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
5616 0 0
2
43331.8 0
0
6 74LS83
105 282 267 0 14 29
0 26 26 27 27 35 34 33 32 26
17 16 15 14 36
0
0 0 4848 0
5 74F83
-18 -60 17 -52
2 U2
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 0 0 0 0
1 U
9323 0 0
2
43331.8 0
0
6 74LS83
105 280 420 0 14 29
0 26 26 27 27 31 30 29 28 26
25 24 23 22 37
0
0 0 4848 0
5 74F83
-18 -60 17 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 0 0 0 0
1 U
317 0 0
2
43331.8 0
0
8 Hex Key~
166 123 82 0 11 12
0 28 29 30 31 0 0 0 0 0
9 57
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
3108 0 0
2
43331.8 0
0
8 Hex Key~
166 74 82 0 11 12
0 32 33 34 35 0 0 0 0 0
13 68
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
4299 0 0
2
43331.8 0
0
45
3 1 2 0 0 8320 0 4 10 0 0 6
856 171
856 168
947 168
947 228
960 228
960 220
2 2 3 0 0 12416 0 5 4 0 0 6
860 334
860 317
872 317
872 225
865 225
865 216
2 1 4 0 0 4224 0 6 4 0 0 4
857 277
857 225
847 225
847 216
1 0 5 0 0 4096 0 5 0 0 14 2
860 370
860 369
1 0 6 0 0 4096 0 6 0 0 6 2
857 313
857 312
3 1 6 0 0 4224 0 7 11 0 0 5
816 312
950 312
950 350
962 350
962 342
2 2 7 0 0 8320 0 9 7 0 0 4
703 407
758 407
758 321
771 321
5 1 8 0 0 4224 0 8 7 0 0 4
679 328
763 328
763 303
771 303
14 1 5 0 0 8192 0 13 9 0 0 4
635 369
659 369
659 407
667 407
4 13 9 0 0 4224 0 8 13 0 0 2
634 342
635 342
3 12 10 0 0 4224 0 8 13 0 0 2
634 333
635 333
2 11 11 0 0 4224 0 8 13 0 0 2
634 324
635 324
1 10 12 0 0 4224 0 8 13 0 0 2
634 315
635 315
14 1 5 0 0 4224 0 13 12 0 0 5
635 369
952 369
952 458
965 458
965 450
1 9 13 0 0 8320 0 1 13 0 0 4
502 324
543 324
543 369
571 369
13 4 14 0 0 4224 0 18 13 0 0 4
314 285
548 285
548 315
571 315
12 3 15 0 0 4224 0 18 13 0 0 4
314 276
553 276
553 306
571 306
11 2 16 0 0 4224 0 18 13 0 0 4
314 267
558 267
558 297
571 297
10 1 17 0 0 4224 0 18 13 0 0 4
314 258
563 258
563 288
571 288
2 8 18 0 0 8320 0 14 13 0 0 4
438 478
548 478
548 351
571 351
2 7 19 0 0 4224 0 15 13 0 0 4
437 440
553 440
553 342
571 342
2 6 20 0 0 4224 0 16 13 0 0 4
436 402
558 402
558 333
571 333
2 5 21 0 0 4224 0 17 13 0 0 4
435 365
563 365
563 324
571 324
13 1 22 0 0 4224 0 19 14 0 0 4
312 438
389 438
389 478
402 478
12 1 23 0 0 4224 0 19 15 0 0 4
312 429
393 429
393 440
401 440
11 1 24 0 0 4224 0 19 16 0 0 4
312 420
387 420
387 402
400 402
10 1 25 0 0 4224 0 19 17 0 0 4
312 411
391 411
391 365
399 365
1 9 26 0 0 8192 0 2 19 0 0 4
184 390
205 390
205 465
248 465
1 9 26 0 0 8192 0 2 18 0 0 4
184 390
212 390
212 313
250 313
1 2 26 0 0 0 0 2 19 0 0 4
184 390
235 390
235 393
248 393
1 1 26 0 0 0 0 2 19 0 0 4
184 390
240 390
240 384
248 384
1 2 26 0 0 8192 0 2 18 0 0 4
184 390
217 390
217 241
250 241
1 1 26 0 0 8320 0 2 18 0 0 4
184 390
222 390
222 232
250 232
1 4 27 0 0 8320 0 3 19 0 0 4
185 228
225 228
225 411
248 411
1 3 27 0 0 0 0 3 19 0 0 4
185 228
230 228
230 402
248 402
1 4 27 0 0 0 0 3 18 0 0 4
185 228
237 228
237 259
250 259
1 3 27 0 0 0 0 3 18 0 0 4
185 228
242 228
242 250
250 250
1 8 28 0 0 4224 0 20 19 0 0 3
132 106
132 447
248 447
2 7 29 0 0 4224 0 20 19 0 0 3
126 106
126 438
248 438
3 6 30 0 0 4224 0 20 19 0 0 3
120 106
120 429
248 429
4 5 31 0 0 4224 0 20 19 0 0 3
114 106
114 420
248 420
1 8 32 0 0 4224 0 21 18 0 0 3
83 106
83 295
250 295
2 7 33 0 0 4224 0 21 18 0 0 3
77 106
77 286
250 286
3 6 34 0 0 8320 0 21 18 0 0 3
71 106
71 277
250 277
4 5 35 0 0 8320 0 21 18 0 0 3
65 106
65 268
250 268
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
501 559 642 583
511 567 631 583
15 XS-3 COMPARATOR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
968 420 1013 444
978 428 1002 444
3 A>B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
966 313 1011 337
976 321 1000 337
3 A=B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
965 189 1010 213
975 197 999 213
3 A<B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
108 19 137 43
118 27 126 43
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
60 20 89 44
70 28 78 44
1 A
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
