CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
110 60 30 120 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
20
13 Logic Switch~
5 292 303 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 514 245 0 1 11
0 8
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
43306.4 0
0
13 Logic Switch~
5 127 438 0 1 11
0 31
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3124 0 0
2
43306.4 1
0
13 Logic Switch~
5 124 243 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
43306.4 2
0
12 Hex Display~
7 744 153 0 18 19
10 4 5 6 7 0 0 0 0 0
0 1 1 1 1 0 1 1 9
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
8157 0 0
2
43306.4 3
0
9 Inverter~
13 416 385 0 2 22
0 10 9
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
5572 0 0
2
43306.4 4
0
5 4030~
219 512 527 0 3 22
0 15 9 11
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U6D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 2 0
1 U
8901 0 0
2
43306.4 5
0
5 4030~
219 513 476 0 3 22
0 16 9 12
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U6C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
7361 0 0
2
43306.4 6
0
5 4030~
219 513 424 0 3 22
0 17 9 13
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U6B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
4747 0 0
2
43306.4 7
0
5 4030~
219 512 370 0 3 22
0 18 9 14
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U6A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
972 0 0
2
43306.4 8
0
6 74LS83
105 627 286 0 14 29
0 8 8 8 8 14 13 12 11 9
7 6 5 4 40
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U5
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
3472 0 0
2
43306.4 9
0
9 Inverter~
13 322 499 0 2 22
0 27 23
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
9998 0 0
2
43306.4 10
0
9 Inverter~
13 322 459 0 2 22
0 28 24
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3536 0 0
2
43306.4 11
0
9 Inverter~
13 322 421 0 2 22
0 29 25
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
4597 0 0
2
43306.4 12
0
9 Inverter~
13 321 384 0 2 22
0 30 26
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3835 0 0
2
43306.4 13
0
6 74LS83
105 397 290 0 14 29
0 22 21 20 19 26 25 24 23 3
18 17 16 15 10
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U3
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
3670 0 0
2
43306.4 14
0
8 Hex Key~
166 142 308 0 11 12
0 32 33 34 35 0 0 0 0 0
9 57
0
0 0 4640 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
5616 0 0
2
43306.4 15
0
8 Hex Key~
166 140 95 0 11 12
0 36 37 38 39 0 0 0 0 0
0 48
0
0 0 4640 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
9323 0 0
2
43306.4 16
0
6 74LS83
105 230 394 0 14 29
0 35 34 33 32 31 31 2 2 31
30 29 28 27 41
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U2
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
317 0 0
2
43306.4 17
0
6 74LS83
105 231 221 0 14 29
0 39 38 37 36 31 31 2 2 31
22 21 20 19 42
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
3108 0 0
2
43306.4 18
0
53
1 8 2 0 0 8320 0 4 19 0 0 4
136 243
175 243
175 421
198 421
1 8 2 0 0 0 0 4 20 0 0 4
136 243
186 243
186 248
199 248
1 9 3 0 0 4224 0 1 16 0 0 4
304 303
342 303
342 335
365 335
13 1 4 0 0 8320 0 11 5 0 0 3
659 304
753 304
753 177
12 2 5 0 0 8320 0 11 5 0 0 3
659 295
747 295
747 177
11 3 6 0 0 8320 0 11 5 0 0 3
659 286
741 286
741 177
10 4 7 0 0 8320 0 11 5 0 0 3
659 277
735 277
735 177
1 4 8 0 0 4096 0 2 11 0 0 4
526 245
572 245
572 277
595 277
1 3 8 0 0 4096 0 2 11 0 0 4
526 245
577 245
577 268
595 268
1 2 8 0 0 4096 0 2 11 0 0 4
526 245
582 245
582 259
595 259
1 1 8 0 0 4224 0 2 11 0 0 4
526 245
587 245
587 250
595 250
2 9 9 0 0 12288 0 6 11 0 0 4
437 385
492 385
492 331
595 331
2 2 9 0 0 8320 0 6 7 0 0 4
437 385
458 385
458 536
496 536
2 2 9 0 0 0 0 6 8 0 0 4
437 385
464 385
464 485
497 485
2 2 9 0 0 0 0 6 9 0 0 4
437 385
469 385
469 433
497 433
2 2 9 0 0 0 0 6 10 0 0 4
437 385
488 385
488 379
496 379
14 1 10 0 0 8320 0 16 6 0 0 6
429 335
441 335
441 400
393 400
393 385
401 385
3 8 11 0 0 8320 0 7 11 0 0 4
545 527
572 527
572 313
595 313
3 7 12 0 0 8320 0 8 11 0 0 4
546 476
577 476
577 304
595 304
3 6 13 0 0 8320 0 9 11 0 0 4
546 424
582 424
582 295
595 295
3 5 14 0 0 8320 0 10 11 0 0 4
545 370
587 370
587 286
595 286
13 1 15 0 0 8320 0 16 7 0 0 4
429 308
473 308
473 518
496 518
12 1 16 0 0 8320 0 16 8 0 0 4
429 299
479 299
479 467
497 467
11 1 17 0 0 8320 0 16 9 0 0 4
429 290
484 290
484 415
497 415
10 1 18 0 0 8320 0 16 10 0 0 4
429 281
488 281
488 361
496 361
13 4 19 0 0 4224 0 20 16 0 0 4
263 239
342 239
342 281
365 281
12 3 20 0 0 4224 0 20 16 0 0 4
263 230
347 230
347 272
365 272
11 2 21 0 0 4224 0 20 16 0 0 4
263 221
352 221
352 263
365 263
10 1 22 0 0 4224 0 20 16 0 0 4
263 212
357 212
357 254
365 254
2 8 23 0 0 8320 0 12 16 0 0 4
343 499
347 499
347 317
365 317
2 7 24 0 0 8320 0 13 16 0 0 4
343 459
347 459
347 308
365 308
2 6 25 0 0 8320 0 14 16 0 0 4
343 421
352 421
352 299
365 299
2 5 26 0 0 8320 0 15 16 0 0 4
342 384
357 384
357 290
365 290
13 1 27 0 0 8320 0 19 12 0 0 4
262 412
289 412
289 499
307 499
12 1 28 0 0 8320 0 19 13 0 0 4
262 403
294 403
294 459
307 459
11 1 29 0 0 4224 0 19 14 0 0 4
262 394
299 394
299 421
307 421
10 1 30 0 0 4224 0 19 15 0 0 4
262 385
298 385
298 384
306 384
1 6 31 0 0 8192 0 3 20 0 0 4
139 438
166 438
166 230
199 230
1 5 31 0 0 8320 0 3 20 0 0 4
139 438
166 438
166 221
199 221
1 9 31 0 0 0 0 3 20 0 0 4
139 438
166 438
166 266
199 266
1 5 31 0 0 0 0 3 19 0 0 4
139 438
170 438
170 394
198 394
1 6 31 0 0 0 0 3 19 0 0 4
139 438
185 438
185 403
198 403
1 9 31 0 0 0 0 3 19 0 0 4
139 438
190 438
190 439
198 439
1 7 2 0 0 0 0 4 19 0 0 4
136 243
180 243
180 412
198 412
1 7 2 0 0 0 0 4 20 0 0 4
136 243
191 243
191 239
199 239
1 4 32 0 0 4224 0 17 19 0 0 3
151 332
151 385
198 385
2 3 33 0 0 8320 0 17 19 0 0 3
145 332
145 376
198 376
3 2 34 0 0 8320 0 17 19 0 0 3
139 332
139 367
198 367
4 1 35 0 0 8320 0 17 19 0 0 3
133 332
133 358
198 358
1 4 36 0 0 4224 0 18 20 0 0 3
149 119
149 212
199 212
2 3 37 0 0 4224 0 18 20 0 0 3
143 119
143 203
199 203
3 2 38 0 0 4224 0 18 20 0 0 3
137 119
137 194
199 194
4 1 39 0 0 8320 0 18 20 0 0 3
131 119
131 185
199 185
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
343 121 528 142
351 128 519 143
21 XS-3 SUBTRACTOR (2'S)
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
