CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
380 70 3 180 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
4
12 Hex Display~
7 506 110 0 18 19
10 2 3 4 5 0 0 0 0 0
0 1 1 1 1 1 1 1 8
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
5130 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 505 195 0 3 22
0 5 3 6
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U2A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
391 0 0
2
5.89855e-315 0
0
7 Pulser~
4 418 335 0 10 12
0 8 9 7 10 0 0 5 5 4
7
0
0 0 4640 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3124 0 0
2
5.89855e-315 0
0
6 74LS93
109 503 273 0 8 17
0 6 6 7 2 5 4 3 2
0
0 0 4832 0
6 74LS93
-21 -35 21 -27
2 U1
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
3421 0 0
2
5.89855e-315 0
0
10
8 1 2 0 0 8320 0 4 1 0 0 5
535 291
564 291
564 157
515 157
515 134
7 2 3 0 0 8320 0 4 1 0 0 5
535 282
559 282
559 152
509 152
509 134
6 3 4 0 0 8320 0 4 1 0 0 5
535 273
554 273
554 147
503 147
503 134
5 4 5 0 0 8320 0 4 1 0 0 5
535 264
549 264
549 142
497 142
497 134
3 2 6 0 0 8320 0 2 4 0 0 4
478 195
452 195
452 273
471 273
3 1 6 0 0 0 0 2 4 0 0 4
478 195
457 195
457 264
471 264
7 2 3 0 0 0 0 4 2 0 0 4
535 282
544 282
544 186
523 186
5 1 5 0 0 0 0 4 2 0 0 4
535 264
539 264
539 204
523 204
8 4 2 0 0 0 0 4 4 0 0 6
535 291
539 291
539 306
452 306
452 291
465 291
3 3 7 0 0 8320 0 3 4 0 0 4
442 326
457 326
457 282
465 282
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 19
436 368 609 392
446 376 598 392
19 DIVIDE BY 9 COUNTER
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
