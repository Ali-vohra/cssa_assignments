CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
14
13 Logic Switch~
5 432 517 0 1 11
0 3
0
0 0 21360 90
2 0V
11 0 25 8
2 V7
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89862e-315 0
0
13 Logic Switch~
5 331 518 0 1 11
0 10
0
0 0 21360 90
2 0V
11 0 25 8
2 V6
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89862e-315 0
0
13 Logic Switch~
5 144 220 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89862e-315 0
0
13 Logic Switch~
5 145 171 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.89862e-315 0
0
13 Logic Switch~
5 147 123 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.89862e-315 0
0
13 Logic Switch~
5 148 81 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
5.89862e-315 0
0
14 Logic Display~
6 901 119 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8901 0 0
2
5.89862e-315 0
0
8 4-In OR~
219 675 140 0 5 22
0 8 7 6 5 4
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U4A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 4 0
1 U
7361 0 0
2
5.89862e-315 0
0
9 4-In AND~
219 522 232 0 5 22
0 11 2 2 9 5
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U3B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 3 0
1 U
4747 0 0
2
5.89862e-315 0
0
9 4-In AND~
219 522 184 0 5 22
0 12 2 2 10 6
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U3A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 3 0
1 U
972 0 0
2
5.89862e-315 0
0
9 4-In AND~
219 522 136 0 5 22
0 13 3 3 9 7
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U2B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 2 0
1 U
3472 0 0
2
5.89862e-315 0
0
9 4-In AND~
219 521 94 0 5 22
0 14 3 3 10 8
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 U2A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 2 0
1 U
9998 0 0
2
5.89862e-315 0
0
9 Inverter~
13 393 465 0 2 22
0 3 2
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U1B
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
3536 0 0
2
5.89862e-315 0
0
9 Inverter~
13 294 464 0 2 22
0 10 9
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U1A
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
4597 0 0
2
5.89862e-315 0
0
27
2 0 2 0 0 4096 0 9 0 0 24 2
498 228
396 228
2 0 2 0 0 0 0 10 0 0 24 2
498 180
396 180
2 0 3 0 0 4096 0 11 0 0 22 2
498 132
433 132
2 0 3 0 0 0 0 12 0 0 22 2
497 90
433 90
5 1 4 0 0 4224 0 8 7 0 0 3
708 140
901 140
901 137
5 4 5 0 0 4224 0 9 8 0 0 4
543 232
633 232
633 154
658 154
5 3 6 0 0 12416 0 10 8 0 0 4
543 184
558 184
558 145
658 145
5 2 7 0 0 4224 0 11 8 0 0 2
543 136
658 136
5 1 8 0 0 4224 0 12 8 0 0 4
542 94
638 94
638 127
658 127
4 0 9 0 0 4096 0 9 0 0 26 2
498 246
297 246
3 0 2 0 0 0 0 9 0 0 24 2
498 237
396 237
4 0 10 0 0 4096 0 10 0 0 23 2
498 198
332 198
3 0 2 0 0 0 0 10 0 0 24 2
498 189
396 189
4 0 9 0 0 0 0 11 0 0 26 2
498 150
297 150
3 0 3 0 0 0 0 11 0 0 22 2
498 141
433 141
4 0 10 0 0 0 0 12 0 0 23 2
497 108
332 108
3 0 3 0 0 0 0 12 0 0 22 2
497 99
433 99
1 1 11 0 0 12416 0 3 9 0 0 4
156 220
171 220
171 219
498 219
1 1 12 0 0 4224 0 4 10 0 0 2
157 171
498 171
1 1 13 0 0 4224 0 5 11 0 0 2
159 123
498 123
1 1 14 0 0 4224 0 6 12 0 0 2
160 81
497 81
0 0 3 0 0 4224 0 0 0 25 0 2
433 492
433 15
0 0 10 0 0 4224 0 0 0 27 0 2
332 490
332 16
2 0 2 0 0 4224 0 13 0 0 0 2
396 447
396 15
1 1 3 0 0 0 0 1 13 0 0 4
433 504
433 491
396 491
396 483
2 0 9 0 0 4224 0 14 0 0 0 2
297 446
297 15
1 1 10 0 0 0 0 2 14 0 0 4
332 505
332 490
297 490
297 482
7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
75 58 112 82
85 66 101 82
2 A3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
73 105 110 129
83 113 99 129
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
72 151 109 175
82 159 98 175
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
73 200 110 224
83 208 99 224
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
427 547 464 571
437 555 453 571
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
323 546 360 570
333 554 349 570
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
932 116 961 140
942 124 950 140
1 D
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
