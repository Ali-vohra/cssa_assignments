CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
210 40 30 170 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
6
13 Logic Switch~
5 398 337 0 1 11
0 7
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89855e-315 0
0
14 Logic Display~
6 852 313 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
391 0 0
2
5.89855e-315 0
0
12 Hex Display~
7 764 152 0 18 19
10 3 4 5 6 0 0 0 0 0
0 1 0 1 1 0 1 1 5
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3124 0 0
2
5.89855e-315 0
0
8 Hex Key~
166 233 152 0 11 12
0 8 9 10 11 0 0 0 0 0
5 53
0
0 0 4640 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3421 0 0
2
5.89855e-315 0
0
8 Hex Key~
166 352 155 0 11 12
0 12 13 14 15 0 0 0 0 0
0 48
0
0 0 4640 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
8157 0 0
2
5.89855e-315 0
0
6 74LS83
105 458 280 0 14 29
0 15 14 13 12 11 10 9 8 7
6 5 4 3 2
0
0 0 4832 0
7 74LS83A
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
5572 0 0
2
5.89855e-315 0
0
14
14 1 2 0 0 4224 0 6 2 0 0 5
490 325
840 325
840 339
852 339
852 331
1 13 3 0 0 8320 0 3 6 0 0 3
773 176
773 298
490 298
2 12 4 0 0 8320 0 3 6 0 0 3
767 176
767 289
490 289
3 11 5 0 0 8320 0 3 6 0 0 3
761 176
761 280
490 280
4 10 6 0 0 8320 0 3 6 0 0 3
755 176
755 271
490 271
1 9 7 0 0 8320 0 1 6 0 0 4
410 337
418 337
418 325
426 325
1 8 8 0 0 8320 0 4 6 0 0 3
242 176
242 307
426 307
2 7 9 0 0 8320 0 4 6 0 0 3
236 176
236 298
426 298
3 6 10 0 0 8320 0 4 6 0 0 3
230 176
230 289
426 289
4 5 11 0 0 8320 0 4 6 0 0 3
224 176
224 280
426 280
1 4 12 0 0 4224 0 5 6 0 0 3
361 179
361 271
426 271
2 3 13 0 0 4224 0 5 6 0 0 3
355 179
355 262
426 262
3 2 14 0 0 8320 0 5 6 0 0 3
349 179
349 253
426 253
4 1 15 0 0 8320 0 5 6 0 0 3
343 179
343 244
426 244
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
429 47 546 71
439 55 535 71
12 BINARY ADDER
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
