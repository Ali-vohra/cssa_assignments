CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
60 10 30 130 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
28
13 Logic Switch~
5 301 286 0 1 11
0 38
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43330.7 0
0
9 2-In AND~
219 779 214 0 3 22
0 4 3 2
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
391 0 0
2
43330.8 0
0
9 Inverter~
13 705 395 0 2 22
0 5 3
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
3124 0 0
2
43330.8 0
0
9 Inverter~
13 705 265 0 2 22
0 6 4
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 2 0
1 U
3421 0 0
2
43330.8 0
0
14 Logic Display~
6 877 193 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8157 0 0
2
43330.8 0
0
14 Logic Display~
6 880 299 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5572 0 0
2
43330.8 0
0
14 Logic Display~
6 876 424 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8901 0 0
2
43330.8 0
0
9 2-In AND~
219 644 335 0 3 22
0 8 7 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
7361 0 0
2
43330.8 0
0
9 2-In AND~
219 573 450 0 3 22
0 10 9 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
4747 0 0
2
43330.8 0
0
9 2-In AND~
219 571 275 0 3 22
0 11 12 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
972 0 0
2
43330.8 0
0
5 4082~
219 573 388 0 5 22
0 17 16 15 14 9
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U5B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 3 0
1 U
3472 0 0
2
43330.8 0
0
5 4082~
219 571 216 0 5 22
0 21 20 19 18 11
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U5A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 3 0
1 U
9998 0 0
2
43330.8 0
0
9 Inverter~
13 494 442 0 2 22
0 5 10
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
3536 0 0
2
43330.8 0
0
9 Inverter~
13 495 286 0 2 22
0 13 12
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
4597 0 0
2
43330.8 0
0
9 Inverter~
13 301 435 0 2 22
0 25 30
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
3835 0 0
2
43330.8 0
0
9 Inverter~
13 301 404 0 2 22
0 24 31
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
3670 0 0
2
43330.8 0
0
9 Inverter~
13 301 372 0 2 22
0 23 32
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
5616 0 0
2
43330.8 0
0
9 Inverter~
13 301 339 0 2 22
0 22 33
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
9323 0 0
2
43330.8 0
0
6 74LS83
105 427 397 0 14 29
0 26 27 28 29 33 32 31 30 13
17 16 15 14 5
0
0 0 4848 0
5 74F83
-18 -60 17 -52
2 U3
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 0 0 0 0
1 U
317 0 0
2
43330.8 0
0
9 Inverter~
13 300 245 0 2 22
0 46 39
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
3108 0 0
2
43330.7 0
0
9 Inverter~
13 300 212 0 2 22
0 45 40
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
4299 0 0
2
43330.7 0
0
9 Inverter~
13 301 177 0 2 22
0 44 41
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
9672 0 0
2
43330.7 0
0
9 Inverter~
13 300 143 0 2 22
0 43 42
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
7876 0 0
2
43330.7 0
0
6 74LS83
105 427 241 0 14 29
0 34 35 36 37 42 41 40 39 38
21 20 19 18 13
0
0 0 4848 0
5 74F83
-18 -60 17 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 0 0 0 0
1 U
6369 0 0
2
43330.7 0
0
8 Hex Key~
166 245 90 0 11 12
0 46 45 44 43 0 0 0 0 0
9 57
0
0 0 4656 0
0
4 KPD4
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
9172 0 0
2
43330.7 0
0
8 Hex Key~
166 205 90 0 11 12
0 25 24 23 22 0 0 0 0 0
6 54
0
0 0 4656 0
0
4 KPD3
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
7100 0 0
2
43330.7 0
0
8 Hex Key~
166 118 89 0 11 12
0 37 36 35 34 0 0 0 0 0
9 57
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
3820 0 0
2
43330.7 0
0
8 Hex Key~
166 76 89 0 11 12
0 29 28 27 26 0 0 0 0 0
7 55
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
7678 0 0
2
43330.7 0
0
49
3 1 2 0 0 4224 0 2 5 0 0 3
800 214
877 214
877 211
2 2 3 0 0 8320 0 3 2 0 0 4
726 395
742 395
742 223
755 223
2 1 4 0 0 8320 0 4 2 0 0 4
726 265
747 265
747 205
755 205
0 1 5 0 0 4096 0 0 3 7 0 3
638 475
638 395
690 395
3 1 6 0 0 8192 0 8 4 0 0 4
665 335
682 335
682 265
690 265
3 1 6 0 0 4224 0 8 6 0 0 3
665 335
880 335
880 317
14 1 5 0 0 12416 0 19 7 0 0 5
459 442
475 442
475 475
876 475
876 442
3 2 7 0 0 8320 0 9 8 0 0 4
594 450
612 450
612 344
620 344
3 1 8 0 0 8320 0 10 8 0 0 4
592 275
612 275
612 326
620 326
5 2 9 0 0 8320 0 11 9 0 0 6
594 388
598 388
598 470
541 470
541 459
549 459
2 1 10 0 0 4224 0 13 9 0 0 4
515 442
541 442
541 441
549 441
14 1 5 0 0 0 0 19 13 0 0 2
459 442
479 442
5 1 11 0 0 8320 0 12 10 0 0 6
592 216
596 216
596 295
534 295
534 266
547 266
2 2 12 0 0 4224 0 14 10 0 0 4
516 286
539 286
539 284
547 284
14 1 13 0 0 4096 0 24 14 0 0 2
459 286
480 286
13 4 14 0 0 4224 0 19 11 0 0 4
459 415
536 415
536 402
549 402
12 3 15 0 0 4224 0 19 11 0 0 4
459 406
541 406
541 393
549 393
11 2 16 0 0 4224 0 19 11 0 0 4
459 397
536 397
536 384
549 384
10 1 17 0 0 4224 0 19 11 0 0 4
459 388
541 388
541 375
549 375
13 4 18 0 0 4224 0 24 12 0 0 4
459 259
524 259
524 230
547 230
12 3 19 0 0 4224 0 24 12 0 0 4
459 250
529 250
529 221
547 221
11 2 20 0 0 4224 0 24 12 0 0 4
459 241
534 241
534 212
547 212
10 1 21 0 0 4224 0 24 12 0 0 4
459 232
539 232
539 203
547 203
4 1 22 0 0 4224 0 26 18 0 0 3
196 114
196 339
286 339
3 1 23 0 0 4224 0 26 17 0 0 3
202 114
202 372
286 372
2 1 24 0 0 4224 0 26 16 0 0 3
208 114
208 404
286 404
1 1 25 0 0 4224 0 26 15 0 0 3
214 114
214 435
286 435
4 1 26 0 0 8320 0 28 19 0 0 5
67 113
67 357
377 357
377 361
395 361
3 2 27 0 0 8320 0 28 19 0 0 5
73 113
73 357
382 357
382 370
395 370
2 3 28 0 0 8320 0 28 19 0 0 5
79 113
79 387
377 387
377 379
395 379
1 4 29 0 0 8320 0 28 19 0 0 3
85 113
85 388
395 388
2 8 30 0 0 4224 0 15 19 0 0 4
322 435
387 435
387 424
395 424
2 7 31 0 0 4224 0 16 19 0 0 4
322 404
387 404
387 415
395 415
2 6 32 0 0 4224 0 17 19 0 0 4
322 372
382 372
382 406
395 406
2 5 33 0 0 4224 0 18 19 0 0 4
322 339
387 339
387 397
395 397
14 9 13 0 0 8320 0 24 19 0 0 6
459 286
463 286
463 457
387 457
387 442
395 442
4 1 34 0 0 8320 0 27 24 0 0 5
109 113
109 197
377 197
377 205
395 205
3 2 35 0 0 8320 0 27 24 0 0 5
115 113
115 227
367 227
367 214
395 214
2 3 36 0 0 8320 0 27 24 0 0 5
121 113
121 227
372 227
372 223
395 223
1 4 37 0 0 8320 0 27 24 0 0 3
127 113
127 232
395 232
1 9 38 0 0 4224 0 1 24 0 0 2
313 286
395 286
2 8 39 0 0 4224 0 20 24 0 0 4
321 245
387 245
387 268
395 268
2 7 40 0 0 4224 0 21 24 0 0 4
321 212
377 212
377 259
395 259
2 6 41 0 0 8320 0 22 24 0 0 4
322 177
382 177
382 250
395 250
2 5 42 0 0 8320 0 23 24 0 0 4
321 143
387 143
387 241
395 241
4 1 43 0 0 8320 0 25 23 0 0 3
236 114
236 143
285 143
3 1 44 0 0 4224 0 25 22 0 0 3
242 114
242 177
286 177
2 1 45 0 0 4224 0 25 21 0 0 3
248 114
248 212
285 212
1 1 46 0 0 4224 0 25 20 0 0 3
254 114
254 245
285 245
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
891 415 934 437
900 422 924 438
3 A>B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
891 289 934 311
900 296 924 312
3 A=B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
891 179 934 201
900 186 924 202
3 A<B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
212 20 241 44
222 28 230 44
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
85 19 114 43
95 27 103 43
1 A
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
