CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
14
13 Logic Switch~
5 738 232 0 1 11
0 2
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 611 266 0 1 11
0 8
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 395 324 0 1 11
0 14
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 145 468 0 1 11
0 23
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 159 255 0 10 11
0 24 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8157 0 0
2
5.89855e-315 0
0
12 Hex Display~
7 886 171 0 18 19
10 3 4 5 6 0 0 0 0 0
0 1 1 1 1 1 1 1 8
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
5572 0 0
2
5.89855e-315 0
0
12 Hex Display~
7 817 173 0 18 19
10 7 2 2 2 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
8901 0 0
2
5.89855e-315 0
0
9 Inverter~
13 589 364 0 2 22
0 7 9
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U5A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
7361 0 0
2
5.89855e-315 0
0
6 74LS83
105 736 310 0 14 29
0 9 8 9 8 13 12 11 10 8
6 5 4 3 33
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U4
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
4747 0 0
2
5.89855e-315 0
0
6 74LS83
105 500 314 0 14 29
0 22 21 20 19 18 17 16 15 14
13 12 11 10 7
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U3
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
972 0 0
2
5.89855e-315 0
0
8 Hex Key~
166 119 342 0 11 12
0 25 26 27 28 0 0 0 0 0
9 57
0
0 0 4640 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3472 0 0
2
5.89855e-315 0
0
8 Hex Key~
166 117 85 0 11 12
0 29 30 31 32 0 0 0 0 0
9 57
0
0 0 4640 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
9998 0 0
2
5.89855e-315 0
0
6 74LS83
105 276 440 0 14 29
0 28 27 26 25 23 23 24 24 23
18 17 16 15 34
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U2
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
3536 0 0
2
5.89855e-315 0
0
6 74LS83
105 274 220 0 14 29
0 32 31 30 29 23 23 24 24 23
22 21 20 19 35
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
4597 0 0
2
5.89855e-315 0
0
45
1 2 2 0 0 4224 0 1 7 0 0 3
750 232
820 232
820 197
1 3 2 0 0 0 0 1 7 0 0 3
750 232
814 232
814 197
1 4 2 0 0 0 0 1 7 0 0 3
750 232
808 232
808 197
13 1 3 0 0 8320 0 9 6 0 0 3
768 328
895 328
895 195
12 2 4 0 0 8320 0 9 6 0 0 3
768 319
889 319
889 195
11 3 5 0 0 4224 0 9 6 0 0 3
768 310
883 310
883 195
10 4 6 0 0 4224 0 9 6 0 0 3
768 301
877 301
877 195
14 1 7 0 0 12416 0 10 7 0 0 5
532 359
570 359
570 205
826 205
826 197
1 9 8 0 0 8320 0 2 9 0 0 4
623 266
676 266
676 355
704 355
1 4 8 0 0 0 0 2 9 0 0 4
623 266
681 266
681 301
704 301
1 2 8 0 0 0 0 2 9 0 0 4
623 266
696 266
696 283
704 283
2 3 9 0 0 4096 0 8 9 0 0 4
610 364
686 364
686 292
704 292
2 1 9 0 0 8320 0 8 9 0 0 4
610 364
691 364
691 274
704 274
14 1 7 0 0 0 0 10 8 0 0 4
532 359
566 359
566 364
574 364
13 8 10 0 0 4224 0 10 9 0 0 4
532 332
696 332
696 337
704 337
12 7 11 0 0 4224 0 10 9 0 0 4
532 323
696 323
696 328
704 328
11 6 12 0 0 4224 0 10 9 0 0 4
532 314
696 314
696 319
704 319
10 5 13 0 0 4224 0 10 9 0 0 4
532 305
696 305
696 310
704 310
1 9 14 0 0 8320 0 3 10 0 0 4
407 324
440 324
440 359
468 359
13 8 15 0 0 4224 0 13 10 0 0 4
308 458
445 458
445 341
468 341
12 7 16 0 0 4224 0 13 10 0 0 4
308 449
450 449
450 332
468 332
11 6 17 0 0 4224 0 13 10 0 0 4
308 440
455 440
455 323
468 323
10 5 18 0 0 4224 0 13 10 0 0 4
308 431
460 431
460 314
468 314
13 4 19 0 0 4224 0 14 10 0 0 4
306 238
445 238
445 305
468 305
12 3 20 0 0 4224 0 14 10 0 0 4
306 229
450 229
450 296
468 296
11 2 21 0 0 4224 0 14 10 0 0 4
306 220
455 220
455 287
468 287
10 1 22 0 0 4224 0 14 10 0 0 4
306 211
460 211
460 278
468 278
1 9 23 0 0 8192 0 4 14 0 0 4
157 468
199 468
199 265
242 265
1 8 24 0 0 8320 0 5 13 0 0 4
171 255
206 255
206 467
244 467
1 7 24 0 0 0 0 5 13 0 0 4
171 255
211 255
211 458
244 458
1 6 23 0 0 8192 0 4 14 0 0 4
157 468
214 468
214 229
242 229
1 5 23 0 0 8320 0 4 14 0 0 4
157 468
219 468
219 220
242 220
1 6 23 0 0 0 0 4 13 0 0 4
157 468
226 468
226 449
244 449
1 5 23 0 0 0 0 4 13 0 0 4
157 468
231 468
231 440
244 440
1 9 23 0 0 0 0 4 13 0 0 4
157 468
236 468
236 485
244 485
1 8 24 0 0 0 0 5 14 0 0 4
171 255
229 255
229 247
242 247
1 7 24 0 0 0 0 5 14 0 0 4
171 255
234 255
234 238
242 238
1 4 25 0 0 8320 0 11 13 0 0 3
128 366
128 431
244 431
2 3 26 0 0 8320 0 11 13 0 0 3
122 366
122 422
244 422
3 2 27 0 0 8320 0 11 13 0 0 3
116 366
116 413
244 413
4 1 28 0 0 8320 0 11 13 0 0 3
110 366
110 404
244 404
1 4 29 0 0 8320 0 12 14 0 0 3
126 109
126 211
242 211
2 3 30 0 0 8320 0 12 14 0 0 3
120 109
120 202
242 202
3 2 31 0 0 8320 0 12 14 0 0 3
114 109
114 193
242 193
4 1 32 0 0 8320 0 12 14 0 0 3
108 109
108 184
242 184
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
453 101 554 125
463 109 543 125
10 XS-3 ADDER
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
