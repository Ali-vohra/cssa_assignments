CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 150 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
24
13 Logic Switch~
5 133 371 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
961 0 0
2
43355 0
0
13 Logic Switch~
5 135 323 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3178 0 0
2
43355 0
0
13 Logic Switch~
5 136 261 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3409 0 0
2
43355 0
0
13 Logic Switch~
5 136 194 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3951 0 0
2
43355 0
0
13 Logic Switch~
5 136 133 0 10 11
0 22 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8885 0 0
2
43355 0
0
13 Logic Switch~
5 137 75 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3780 0 0
2
43355 0
0
14 Logic Display~
6 928 783 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L16
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9265 0 0
2
43355 0
0
14 Logic Display~
6 925 734 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L15
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9442 0 0
2
43355 0
0
14 Logic Display~
6 924 681 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L14
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9424 0 0
2
43355 0
0
14 Logic Display~
6 922 629 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L13
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9968 0 0
2
43355 0
0
14 Logic Display~
6 920 580 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9281 0 0
2
43355 0
0
14 Logic Display~
6 919 529 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8464 0 0
2
43355 0
0
14 Logic Display~
6 917 478 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7168 0 0
2
43355 0
0
14 Logic Display~
6 915 430 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3171 0 0
2
43355 0
0
14 Logic Display~
6 913 378 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4139 0 0
2
43355 0
0
14 Logic Display~
6 912 322 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6435 0 0
2
43355 0
0
14 Logic Display~
6 911 274 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5283 0 0
2
43355 0
0
14 Logic Display~
6 909 223 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6874 0 0
2
43355 0
0
14 Logic Display~
6 908 172 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5305 0 0
2
43355 0
0
14 Logic Display~
6 907 122 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
34 0 0
2
43355 0
0
14 Logic Display~
6 907 72 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
969 0 0
2
43355 0
0
14 Logic Display~
6 907 24 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8402 0 0
2
43355 0
0
7 74LS138
19 439 311 0 14 29
0 22 21 20 23 18 18 17 16 15
14 13 12 11 10
0
0 0 5104 0
7 74LS138
-25 -61 24 -53
2 U2
-7 -71 7 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 0 0 0 0
1 U
3751 0 0
2
43355 0
0
7 74LS138
19 440 76 0 14 29
0 22 21 20 19 23 23 9 8 7
6 5 4 3 2
0
0 0 5104 0
7 74LS138
-25 -61 24 -53
2 U1
-7 -71 7 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 0 0 0 0
1 U
4292 0 0
2
43355 0
0
28
14 1 2 0 0 8320 0 24 7 0 0 4
478 112
801 112
801 801
928 801
13 1 3 0 0 8320 0 24 8 0 0 4
478 103
810 103
810 752
925 752
12 1 4 0 0 8320 0 24 9 0 0 4
478 94
819 94
819 699
924 699
11 1 5 0 0 8320 0 24 10 0 0 4
478 85
827 85
827 647
922 647
10 1 6 0 0 8320 0 24 11 0 0 4
478 76
836 76
836 598
920 598
9 1 7 0 0 8320 0 24 12 0 0 4
478 67
843 67
843 547
919 547
8 1 8 0 0 8320 0 24 13 0 0 4
478 58
850 58
850 496
917 496
7 1 9 0 0 8320 0 24 14 0 0 4
478 49
857 49
857 448
915 448
14 1 10 0 0 4224 0 23 15 0 0 5
477 347
876 347
876 404
913 404
913 396
13 1 11 0 0 4224 0 23 16 0 0 5
477 338
880 338
880 349
912 349
912 340
12 1 12 0 0 4224 0 23 17 0 0 5
477 329
875 329
875 299
911 299
911 292
11 1 13 0 0 4224 0 23 18 0 0 5
477 320
880 320
880 249
909 249
909 241
10 1 14 0 0 4224 0 23 19 0 0 5
477 311
863 311
863 198
908 198
908 190
9 1 15 0 0 4224 0 23 20 0 0 5
477 302
867 302
867 148
907 148
907 140
8 1 16 0 0 4224 0 23 21 0 0 5
477 293
871 293
871 99
907 99
907 90
7 1 17 0 0 4224 0 23 22 0 0 5
477 284
876 284
876 51
907 51
907 42
1 6 18 0 0 4096 0 1 23 0 0 4
145 371
388 371
388 347
401 347
1 5 18 0 0 4224 0 1 23 0 0 4
145 371
393 371
393 338
401 338
1 4 19 0 0 4224 0 2 24 0 0 4
147 323
394 323
394 94
408 94
1 3 20 0 0 4224 0 3 23 0 0 4
148 261
387 261
387 302
407 302
1 2 21 0 0 4224 0 4 23 0 0 4
148 194
382 194
382 293
407 293
1 1 22 0 0 4224 0 5 23 0 0 4
148 133
387 133
387 284
407 284
1 3 20 0 0 0 0 3 24 0 0 4
148 261
362 261
362 67
408 67
1 2 21 0 0 0 0 4 24 0 0 4
148 194
367 194
367 58
408 58
1 1 22 0 0 0 0 5 24 0 0 4
148 133
372 133
372 49
408 49
1 4 23 0 0 8320 0 6 23 0 0 4
149 75
377 75
377 329
407 329
1 6 23 0 0 0 0 6 24 0 0 4
149 75
382 75
382 112
402 112
1 5 23 0 0 0 0 6 24 0 0 4
149 75
387 75
387 103
402 103
20
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
938 769 975 793
948 777 964 793
2 D0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
937 719 974 743
947 727 963 743
2 D1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
935 666 972 690
945 674 961 690
2 D2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
933 614 970 638
943 622 959 638
2 D3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
931 565 968 589
941 573 957 589
2 D4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
930 515 967 539
940 523 956 539
2 D5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
930 464 967 488
940 472 956 488
2 D6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
928 414 965 438
938 422 954 438
2 D7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
926 364 963 388
936 372 952 388
2 D8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
924 309 961 333
934 317 950 333
2 D9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
922 261 967 285
932 269 956 285
3 D10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
922 210 967 234
932 218 956 234
3 D11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
920 159 965 183
930 167 954 183
3 D12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
918 109 963 133
928 117 952 133
3 D13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
917 58 962 82
927 66 951 82
3 D14
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
916 9 961 33
926 17 950 33
3 D15
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
74 237 111 261
84 245 100 261
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
73 172 110 196
83 180 99 196
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
73 108 110 132
83 116 99 132
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
74 51 111 75
84 59 100 75
2 A3
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
