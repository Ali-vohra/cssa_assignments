CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 90 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
36
13 Logic Switch~
5 105 814 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V11
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43382.9 0
0
13 Logic Switch~
5 106 766 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V10
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
43382.9 0
0
13 Logic Switch~
5 105 715 0 1 11
0 31
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
43382.9 0
0
13 Logic Switch~
5 102 605 0 1 11
0 34
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3421 0 0
2
43382.9 0
0
13 Logic Switch~
5 101 548 0 10 11
0 30 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8157 0 0
2
43382.9 0
0
13 Logic Switch~
5 97 432 0 1 11
0 26
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5572 0 0
2
43382.9 0
0
13 Logic Switch~
5 98 382 0 10 11
0 22 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8901 0 0
2
43382.9 0
0
13 Logic Switch~
5 95 278 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7361 0 0
2
43382.9 0
0
13 Logic Switch~
5 96 230 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4747 0 0
2
43382.9 0
0
13 Logic Switch~
5 93 137 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
972 0 0
2
43382.9 0
0
13 Logic Switch~
5 93 94 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3472 0 0
2
43382.9 0
0
14 Logic Display~
6 1147 1194 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9998 0 0
2
43382.9 0
0
14 Logic Display~
6 899 1195 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3536 0 0
2
43382.9 0
0
9 2-In AND~
219 873 883 0 3 22
0 9 10 12
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U6D
-12 -6 9 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
4597 0 0
2
43382.9 2
0
9 2-In AND~
219 918 884 0 3 22
0 7 8 11
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U6C
-12 -6 9 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
3835 0 0
2
43382.9 1
0
8 2-In OR~
219 890 957 0 3 22
0 11 12 6
0
0 0 624 270
6 74LS32
-21 -24 21 -16
3 U3D
-7 -1 14 7
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
3670 0 0
2
43382.9 0
0
14 Logic Display~
6 687 1199 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5616 0 0
2
43382.9 0
0
9 2-In AND~
219 664 882 0 3 22
0 18 10 20
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U6B
-12 -6 9 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
9323 0 0
2
43382.9 2
0
9 2-In AND~
219 709 883 0 3 22
0 17 8 19
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U6A
-12 -6 9 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
317 0 0
2
43382.9 1
0
8 2-In OR~
219 681 956 0 3 22
0 19 20 16
0
0 0 624 270
6 74LS32
-21 -24 21 -16
3 U3C
-7 -1 14 7
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
3108 0 0
2
43382.9 0
0
14 Logic Display~
6 482 1204 0 1 2
10 21
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4299 0 0
2
43382.9 0
0
9 2-In AND~
219 458 880 0 3 22
0 26 10 28
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U2D
-12 -6 9 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
9672 0 0
2
43382.9 2
0
9 2-In AND~
219 503 881 0 3 22
0 25 8 27
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U2C
-12 -6 9 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
7876 0 0
2
43382.9 1
0
8 2-In OR~
219 475 954 0 3 22
0 27 28 24
0
0 0 624 270
6 74LS32
-21 -24 21 -16
3 U3B
-7 -1 14 7
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
6369 0 0
2
43382.9 0
0
14 Logic Display~
6 265 1208 0 1 2
10 29
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9172 0 0
2
43382.9 0
0
8 2-In OR~
219 260 952 0 3 22
0 35 36 32
0
0 0 624 270
6 74LS32
-21 -24 21 -16
3 U3A
-7 -1 14 7
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
7100 0 0
2
43382.9 0
0
9 2-In AND~
219 288 879 0 3 22
0 33 8 35
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U2B
-12 -6 9 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3820 0 0
2
43382.9 0
0
9 2-In AND~
219 243 878 0 3 22
0 34 10 36
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U2A
-12 -6 9 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
7678 0 0
2
43382.9 0
0
9 Inverter~
13 158 636 0 2 22
0 34 33
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
961 0 0
2
43382.9 0
0
9 Inverter~
13 154 462 0 2 22
0 26 25
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3178 0 0
2
43382.9 0
0
9 Inverter~
13 154 310 0 2 22
0 18 17
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
3409 0 0
2
43382.9 0
0
9 Inverter~
13 152 167 0 2 22
0 9 7
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3951 0 0
2
43382.9 0
0
2 FA
94 264 1049 0 5 11
0 30 32 31 23 29
2 FA
1 0 688 0
0
2 U4
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
8885 0 0
2
43334.9 0
0
2 FA
94 481 1049 0 5 11
0 22 24 23 15 21
2 FA
2 0 688 0
0
2 U5
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
3780 0 0
2
43334.9 0
0
2 FA
94 686 1049 0 5 11
0 14 16 15 5 13
2 FA
3 0 688 0
0
2 U7
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
9265 0 0
2
43334.9 0
0
2 FA
94 897 1049 0 5 11
0 4 6 5 2 3
2 FA
4 0 688 0
0
2 U8
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
9442 0 0
2
43334.9 0
0
60
4 1 2 0 0 8320 0 36 12 0 0 5
930 1067
1088 1067
1088 1237
1147 1237
1147 1212
5 1 3 0 0 12416 0 36 13 0 0 7
930 1049
975 1049
975 1125
808 1125
808 1237
899 1237
899 1213
1 0 4 0 0 8320 0 36 0 0 60 3
864 1049
817 1049
817 94
4 3 5 0 0 4224 0 35 36 0 0 2
719 1067
864 1067
3 2 6 0 0 8320 0 16 36 0 0 5
893 987
893 1003
808 1003
808 1058
864 1058
1 0 7 0 0 4096 0 15 0 0 57 2
925 862
925 167
2 0 8 0 0 4096 0 15 0 0 43 2
907 862
907 766
1 0 9 0 0 4096 0 14 0 0 59 2
880 861
880 137
2 0 10 0 0 4096 0 14 0 0 42 2
862 861
862 814
3 1 11 0 0 4240 0 15 16 0 0 4
916 907
916 926
902 926
902 941
3 2 12 0 0 4240 0 14 16 0 0 4
871 906
871 926
884 926
884 941
5 1 13 0 0 12416 0 35 17 0 0 7
719 1049
749 1049
749 1124
600 1124
600 1236
687 1236
687 1217
1 0 14 0 0 8192 0 35 0 0 56 3
653 1049
608 1049
608 230
4 3 15 0 0 4224 0 34 35 0 0 2
514 1067
653 1067
3 2 16 0 0 8320 0 20 35 0 0 5
684 986
684 1003
600 1003
600 1058
653 1058
1 0 17 0 0 4096 0 19 0 0 53 2
716 861
716 310
2 0 8 0 0 0 0 19 0 0 43 2
698 861
698 766
1 0 18 0 0 4096 0 18 0 0 55 2
671 860
671 278
2 0 10 0 0 0 0 18 0 0 42 2
653 860
653 814
3 1 19 0 0 4224 0 19 20 0 0 4
707 906
707 925
693 925
693 940
3 2 20 0 0 4224 0 18 20 0 0 4
662 905
662 925
675 925
675 940
5 1 21 0 0 12416 0 34 21 0 0 7
514 1049
555 1049
555 1124
399 1124
399 1236
482 1236
482 1222
1 0 22 0 0 8192 0 34 0 0 52 3
448 1049
407 1049
407 382
3 4 23 0 0 4224 0 34 33 0 0 2
448 1067
297 1067
3 2 24 0 0 8320 0 24 34 0 0 5
478 984
478 1002
399 1002
399 1058
448 1058
1 0 25 0 0 4096 0 23 0 0 49 2
510 859
510 462
2 0 8 0 0 0 0 23 0 0 43 2
492 859
492 766
1 0 26 0 0 4096 0 22 0 0 51 2
465 858
465 432
2 0 10 0 0 0 0 22 0 0 42 2
447 858
447 814
3 1 27 0 0 4224 0 23 24 0 0 4
501 904
501 923
487 923
487 938
3 2 28 0 0 4224 0 22 24 0 0 4
456 903
456 923
469 923
469 938
5 1 29 0 0 12416 0 33 25 0 0 7
297 1049
330 1049
330 1124
215 1124
215 1236
265 1236
265 1226
1 0 30 0 0 8192 0 33 0 0 48 3
231 1049
214 1049
214 548
3 0 31 0 0 8192 0 33 0 0 44 3
231 1067
205 1067
205 715
3 2 32 0 0 8320 0 26 33 0 0 5
263 982
263 1004
197 1004
197 1058
231 1058
1 0 33 0 0 4096 0 27 0 0 45 2
295 857
295 636
2 0 8 0 0 0 0 27 0 0 43 2
277 857
277 766
1 0 34 0 0 4096 0 28 0 0 47 2
250 856
250 605
2 0 10 0 0 0 0 28 0 0 42 2
232 856
232 814
3 1 35 0 0 4224 0 27 26 0 0 4
286 902
286 921
272 921
272 936
3 2 36 0 0 4224 0 28 26 0 0 4
241 901
241 921
254 921
254 936
1 0 10 0 0 4224 0 1 0 0 0 2
117 814
1009 814
1 0 8 0 0 4224 0 2 0 0 0 2
118 766
1008 766
1 0 31 0 0 4224 0 3 0 0 0 2
117 715
1008 715
2 0 33 0 0 4224 0 29 0 0 0 2
179 636
1008 636
1 1 34 0 0 0 0 4 29 0 0 4
114 605
135 605
135 636
143 636
1 0 34 0 0 4224 0 4 0 0 0 2
114 605
1009 605
1 0 30 0 0 4224 0 5 0 0 0 2
113 548
1009 548
2 0 25 0 0 4224 0 30 0 0 0 2
175 462
1009 462
1 1 26 0 0 0 0 6 30 0 0 4
109 432
131 432
131 462
139 462
1 0 26 0 0 4224 0 6 0 0 0 2
109 432
1010 432
1 0 22 0 0 4224 0 7 0 0 0 2
110 382
1010 382
2 0 17 0 0 4224 0 31 0 0 0 2
175 310
1011 310
1 1 18 0 0 0 0 8 31 0 0 4
107 278
131 278
131 310
139 310
1 0 18 0 0 4224 0 8 0 0 0 2
107 278
1011 278
1 0 14 0 0 4224 0 9 0 0 0 2
108 230
1012 230
2 0 7 0 0 4224 0 32 0 0 0 2
173 167
1010 167
1 1 9 0 0 0 0 10 32 0 0 4
105 137
129 137
129 167
137 167
1 0 9 0 0 4224 0 10 0 0 0 2
105 137
1011 137
1 0 4 0 0 0 0 11 0 0 0 2
105 94
1011 94
16
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1123 1247 1176 1271
1133 1255 1165 1271
4 Cout
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
883 1253 920 1277
893 1261 909 1277
2 F3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
670 1255 707 1279
680 1263 696 1279
2 F2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
464 1257 501 1281
474 1265 490 1281
2 F1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
246 1261 283 1285
256 1269 272 1285
2 F0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
35 792 72 816
45 800 61 816
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
37 746 74 770
47 754 63 770
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
37 693 82 717
47 701 71 717
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
39 582 76 606
49 590 65 606
2 B0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
39 525 76 549
49 533 65 549
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
33 411 70 435
43 419 59 435
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
35 361 72 385
45 369 61 385
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
36 257 73 281
46 265 62 281
2 B2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
36 211 73 235
46 219 62 235
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
36 115 73 139
46 123 62 139
2 B3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
37 72 74 96
47 80 63 96
2 A3
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
