CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 31 432 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43353.9 0
0
13 Logic Switch~
5 28 488 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
43353.9 0
0
12 Hex Display~
7 494 42 0 16 19
10 3 4 5 6 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3124 0 0
2
43353.9 0
0
12 Hex Display~
7 444 43 0 16 19
10 2 32 33 34 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 0 0 0 0
4 DISP
3421 0 0
2
43353.9 0
0
6 74LS93
109 125 479 0 8 17
0 7 7 19 15 18 17 16 15
0
0 0 4848 0
6 74LS93
-21 -35 21 -27
2 U5
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 0 0 0 0
1 U
8157 0 0
2
43353.9 0
0
8 Hex Key~
166 118 46 0 11 12
0 11 12 13 14 0 0 0 0 0
0 48
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
5572 0 0
2
43353.9 0
0
2 FA
94 302 111 0 5 11
0 14 18 8 2 6
2 FA
1 0 688 0
0
2 U1
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
8901 0 0
2
43334.9 0
0
2 FA
94 302 195 0 5 11
0 13 17 9 8 5
2 FA
2 0 688 0
0
2 U2
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
7361 0 0
2
43334.9 0
0
2 FA
94 302 282 0 5 11
0 12 16 10 9 4
2 FA
3 0 688 0
0
2 U3
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
4747 0 0
2
43334.9 0
0
2 FA
94 302 369 0 5 11
0 11 15 7 10 3
2 FA
4 0 688 0
0
2 U4
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
972 0 0
2
43334.9 0
0
21
4 1 2 0 0 4224 0 7 4 0 0 3
335 129
453 129
453 67
5 1 3 0 0 8320 0 10 3 0 0 3
335 369
503 369
503 66
5 2 4 0 0 8320 0 9 3 0 0 3
335 282
497 282
497 66
5 3 5 0 0 4224 0 8 3 0 0 3
335 195
491 195
491 66
5 4 6 0 0 4224 0 7 3 0 0 3
335 111
485 111
485 66
1 3 7 0 0 4224 0 1 10 0 0 4
43 432
241 432
241 387
269 387
4 3 8 0 0 12416 0 8 7 0 0 5
335 213
353 213
353 156
269 156
269 129
4 3 9 0 0 12416 0 9 8 0 0 5
335 300
353 300
353 242
269 242
269 213
4 3 10 0 0 12416 0 10 9 0 0 5
335 387
353 387
353 329
269 329
269 300
1 1 11 0 0 4224 0 6 10 0 0 3
127 70
127 369
269 369
2 1 12 0 0 4224 0 6 9 0 0 3
121 70
121 282
269 282
3 1 13 0 0 8320 0 6 8 0 0 3
115 70
115 195
269 195
4 1 14 0 0 8320 0 6 7 0 0 3
109 70
109 111
269 111
8 2 15 0 0 8320 0 5 10 0 0 4
157 497
246 497
246 378
269 378
7 2 16 0 0 8320 0 5 9 0 0 4
157 488
251 488
251 291
269 291
6 2 17 0 0 8320 0 5 8 0 0 4
157 479
256 479
256 204
269 204
5 2 18 0 0 8320 0 5 7 0 0 4
157 470
261 470
261 120
269 120
4 8 15 0 0 0 0 5 5 0 0 6
87 497
83 497
83 512
165 512
165 497
157 497
1 2 7 0 0 0 0 1 5 0 0 4
43 432
74 432
74 479
93 479
1 1 7 0 0 0 0 1 5 0 0 4
43 432
79 432
79 470
93 470
1 3 19 0 0 4224 0 2 5 0 0 2
40 488
87 488
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
