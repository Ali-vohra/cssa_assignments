CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
50 50 30 110 9
0 70 1024 728
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 E:\CM60S\BOM.DAT
0 7
0 70 1024 728
143654930 0
0
6 Title:
5 Name:
0
0
0
14
13 Logic Switch~
5 268 281 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 104 203 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 104 157 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 105 115 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6153 0 0
0
0
14 Logic Display~
6 906 290 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5394 0 0
0
0
14 Logic Display~
6 906 340 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7734 0 0
0
0
9 2-In AND~
219 197 179 0 3 22
0 7 9 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
9914 0 0
0
0
14 Logic Display~
6 907 389 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3747 0 0
0
0
9 2-In AND~
219 195 126 0 3 22
0 7 10 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3549 0 0
0
0
6 74LS83
105 390 117 0 14 29
0 2 7 2 9 2 8 6 12 2
3 4 5 11 13
0
0 0 13040 0
7 74LS83A
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
7931 0 0
0
0
9 2-In AND~
219 194 75 0 3 22
0 9 10 12
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
9325 0 0
0
0
14 Logic Display~
6 908 442 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8903 0 0
0
0
14 Logic Display~
6 908 495 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 0 0 0 0
1 L
3834 0 0
0
0
14 Logic Display~
6 909 548 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3363 0 0
0
0
20
1 1 2 0 0 8320 0 1 10 0 0 4
280 281
350 281
350 81
358 81
1 3 2 0 0 0 0 1 10 0 0 4
280 281
350 281
350 99
358 99
1 5 2 0 0 0 0 1 10 0 0 4
280 281
350 281
350 117
358 117
1 9 2 0 0 128 0 1 10 0 0 6
280 281
292 281
292 99
350 99
350 162
358 162
10 1 3 0 0 4224 0 10 5 0 0 5
422 108
893 108
893 316
906 316
906 308
11 1 4 0 0 4224 0 10 6 0 0 5
422 117
893 117
893 366
906 366
906 358
12 1 5 0 0 4224 0 10 8 0 0 5
422 126
894 126
894 415
907 415
907 407
3 7 6 0 0 4224 0 9 10 0 0 4
216 126
350 126
350 135
358 135
1 2 7 0 0 12416 0 4 10 0 0 6
117 115
166 115
166 55
350 55
350 90
358 90
3 6 8 0 0 4224 0 7 10 0 0 4
218 179
350 179
350 126
358 126
1 2 9 0 0 4096 0 3 7 0 0 4
116 157
165 157
165 188
173 188
1 1 7 0 0 0 0 4 7 0 0 4
117 115
165 115
165 170
173 170
1 2 10 0 0 8192 0 2 9 0 0 4
116 203
163 203
163 135
171 135
1 1 7 0 0 0 0 4 9 0 0 4
117 115
163 115
163 117
171 117
13 1 11 0 0 4224 0 10 12 0 0 5
422 135
895 135
895 468
908 468
908 460
1 4 9 0 0 4224 0 3 10 0 0 4
116 157
350 157
350 108
358 108
3 8 12 0 0 4224 0 11 10 0 0 4
215 75
350 75
350 144
358 144
1 2 10 0 0 8192 0 2 11 0 0 4
116 203
162 203
162 84
170 84
1 1 9 0 0 0 0 3 11 0 0 4
116 157
162 157
162 66
170 66
1 1 10 0 0 4224 0 2 14 0 0 5
116 203
896 203
896 574
909 574
909 566
9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
911 279 935 303
921 287 937 303
2 S5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
910 330 934 354
920 338 936 354
2 S4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
912 379 936 403
922 387 938 403
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
915 431 939 455
925 439 941 455
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
913 484 937 508
923 492 939 508
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
913 539 937 563
923 547 939 563
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
55 181 79 205
65 189 81 205
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
55 134 79 158
65 142 81 158
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
56 86 80 110
66 94 82 110
2 A2
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
