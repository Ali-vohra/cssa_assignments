CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
40 10 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
15
13 Logic Switch~
5 148 462 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6118 0 0
2
43355 0
0
13 Logic Switch~
5 149 394 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
34 0 0
2
43355 0
0
13 Logic Switch~
5 149 326 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6357 0 0
2
43355 0
0
13 Logic Switch~
5 148 257 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
319 0 0
2
43355 0
0
13 Logic Switch~
5 148 196 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3976 0 0
2
43355 0
0
14 Logic Display~
6 877 506 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7634 0 0
2
43355 0
0
14 Logic Display~
6 877 444 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
523 0 0
2
43355 0
0
14 Logic Display~
6 876 376 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6748 0 0
2
43355 0
0
14 Logic Display~
6 874 317 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6901 0 0
2
43355 0
0
14 Logic Display~
6 874 257 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
842 0 0
2
43355 0
0
14 Logic Display~
6 872 197 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3277 0 0
2
43355 0
0
14 Logic Display~
6 872 142 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4212 0 0
2
43355 0
0
14 Logic Display~
6 872 81 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4720 0 0
2
43355 0
0
8 2-4 DEC~
94 488 134 0 8 17
0 11 10 14 13 2 3 4 5
8 2-4 DEC~
1 0 816 0
7 2-4 DEC
-22 -92 27 -84
2 U1
-3 -77 11 -69
0
0
0
0
0
0
17

0 1 2 7 8 11 12 13 14 1
2 7 8 11 12 13 14 0
0 0 0 0 1 0 0 0
1 U
5551 0 0
2
43355 0
0
8 2-4 DEC~
94 487 380 0 8 17
0 11 10 12 14 6 7 8 9
8 2-4 DEC~
2 0 816 0
7 2-4 DEC
-23 -88 26 -80
2 U2
-3 -77 11 -69
0
0
0
0
0
0
17

0 1 2 7 8 11 12 13 14 1
2 7 8 11 12 13 14 0
0 0 0 0 1 0 0 0
1 U
6986 0 0
2
43355 0
0
16
5 1 2 0 0 8320 0 14 6 0 0 4
538 161
786 161
786 524
877 524
6 1 3 0 0 8320 0 14 7 0 0 5
538 147
790 147
790 469
877 469
877 462
7 1 4 0 0 8320 0 14 8 0 0 5
538 134
795 134
795 412
876 412
876 394
8 1 5 0 0 4224 0 14 9 0 0 5
538 121
800 121
800 347
874 347
874 335
5 1 6 0 0 4224 0 15 10 0 0 4
537 407
806 407
806 275
874 275
6 1 7 0 0 4224 0 15 11 0 0 5
537 393
810 393
810 223
872 223
872 215
7 1 8 0 0 4224 0 15 12 0 0 5
537 380
815 380
815 163
872 163
872 160
8 1 9 0 0 4224 0 15 13 0 0 5
537 367
820 367
820 105
872 105
872 99
1 2 10 0 0 4224 0 3 15 0 0 4
161 326
422 326
422 353
445 353
1 1 11 0 0 4224 0 4 15 0 0 4
160 257
437 257
437 340
445 340
1 2 10 0 0 0 0 3 14 0 0 4
161 326
418 326
418 107
446 107
1 1 11 0 0 0 0 4 14 0 0 4
160 257
423 257
423 94
446 94
1 3 12 0 0 4224 0 1 15 0 0 4
160 462
437 462
437 420
445 420
1 4 13 0 0 4224 0 2 14 0 0 4
161 394
428 394
428 188
446 188
1 4 14 0 0 4096 0 5 15 0 0 4
160 196
432 196
432 434
445 434
1 3 14 0 0 4224 0 5 14 0 0 4
160 196
438 196
438 174
446 174
11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
884 490 921 514
894 498 910 514
2 D0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
885 429 922 453
895 437 911 453
2 D1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
884 361 921 385
894 369 910 385
2 D2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
884 303 921 327
894 311 910 327
2 D3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
885 241 922 265
895 249 911 265
2 D4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
882 183 919 207
892 191 908 207
2 D5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
882 127 919 151
892 135 908 151
2 D6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
883 67 920 91
893 75 909 91
2 D7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
83 305 120 329
93 313 109 329
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
77 242 114 266
87 250 103 266
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
75 177 112 201
85 185 101 201
2 A2
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
