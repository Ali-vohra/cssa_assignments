CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
10 0 30 80 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
21
13 Logic Switch~
5 159 574 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43354 0
0
13 Logic Switch~
5 30 375 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
43354 0
0
13 Logic Switch~
5 116 575 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3124 0 0
2
43354 0
0
13 Logic Switch~
5 31 432 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.89861e-315 0
0
13 Logic Switch~
5 28 488 0 1 11
0 33
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.89861e-315 0
0
9 Inverter~
13 248 470 0 2 22
0 19 20
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U10E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
5572 0 0
2
43354 0
0
9 Inverter~
13 247 686 0 2 22
0 16 13
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U10D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
8901 0 0
2
43354 0
0
9 Inverter~
13 246 611 0 2 22
0 17 14
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U10C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
7361 0 0
2
43354 0
0
9 Inverter~
13 248 537 0 2 22
0 18 15
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 U10B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
4747 0 0
2
43354 0
0
12 Hex Display~
7 494 42 0 16 19
10 22 23 24 25 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
972 0 0
2
5.89861e-315 0
0
12 Hex Display~
7 444 43 0 16 19
10 21 59 60 61 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
3472 0 0
2
5.89861e-315 0
0
6 74LS93
109 125 479 0 8 17
0 7 7 33 16 19 18 17 16
0
0 0 4848 0
6 74LS93
-21 -35 21 -27
2 U5
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
9998 0 0
2
5.89861e-315 0
0
8 Hex Key~
166 118 46 0 11 12
0 29 30 31 32 0 0 0 0 0
0 48
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3536 0 0
2
5.89861e-315 0
0
2 FA
94 302 111 0 5 11
0 32 6 26 21 25
2 FA
1 0 688 0
0
2 U1
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 1 0 0 0
1 U
4597 0 0
2
5.89859e-315 0
0
2 FA
94 302 195 0 5 11
0 31 5 27 26 24
2 FA
2 0 688 0
0
2 U2
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 1 0 0 0
1 U
3835 0 0
2
5.89859e-315 0
0
2 FA
94 302 282 0 5 11
0 30 4 28 27 23
2 FA
3 0 688 0
0
2 U3
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 1 0 0 0
1 U
3670 0 0
2
5.89859e-315 0
0
2 FA
94 302 369 0 5 11
0 29 3 8 28 22
2 FA
4 0 688 0
0
2 U4
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 1 0 0 0
1 U
5616 0 0
2
5.89859e-315 0
0
2 FA
94 302 470 0 5 11
0 20 2 9 46 6
2 FA
9 0 688 0
0
2 U6
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
9323 0 0
2
43334.9 0
0
2 FA
94 301 537 0 5 11
0 15 2 10 9 5
2 FA
10 0 688 0
0
2 U7
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
317 0 0
2
43334.9 0
0
2 FA
94 299 611 0 5 11
0 14 2 11 10 4
2 FA
11 0 688 0
0
2 U8
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
3108 0 0
2
43334.9 0
0
2 FA
94 298 686 0 5 11
0 13 12 8 11 3
2 FA
12 0 688 0
0
2 U9
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
4299 0 0
2
43334.9 0
0
37
1 2 2 0 0 8192 0 1 20 0 0 3
171 574
171 620
266 620
1 2 2 0 0 8192 0 1 19 0 0 3
171 574
171 546
268 546
1 2 2 0 0 8320 0 1 18 0 0 3
171 574
171 479
269 479
5 2 3 0 0 8320 0 21 17 0 0 6
331 686
359 686
359 345
261 345
261 378
269 378
5 2 4 0 0 8320 0 20 16 0 0 6
332 611
349 611
349 258
261 258
261 291
269 291
5 2 5 0 0 8320 0 19 15 0 0 6
334 537
344 537
344 227
261 227
261 204
269 204
5 2 6 0 0 8320 0 18 14 0 0 6
335 470
339 470
339 87
261 87
261 120
269 120
1 1 7 0 0 8192 0 2 12 0 0 4
42 375
74 375
74 470
93 470
1 2 7 0 0 8320 0 2 12 0 0 4
42 375
79 375
79 479
93 479
1 3 8 0 0 4224 0 4 21 0 0 3
43 432
43 704
265 704
4 3 9 0 0 12416 0 19 18 0 0 6
334 555
339 555
339 502
261 502
261 488
269 488
4 3 10 0 0 12416 0 20 19 0 0 6
332 629
338 629
338 569
260 569
260 555
268 555
4 3 11 0 0 12416 0 21 20 0 0 6
331 704
336 704
336 643
258 643
258 629
266 629
1 2 12 0 0 8320 0 3 21 0 0 3
128 575
128 695
265 695
1 2 13 0 0 4224 0 21 7 0 0 2
265 686
268 686
1 2 14 0 0 4224 0 20 8 0 0 2
266 611
267 611
1 2 15 0 0 4224 0 19 9 0 0 2
268 537
269 537
8 1 16 0 0 8320 0 12 7 0 0 4
157 497
214 497
214 686
232 686
7 1 17 0 0 8320 0 12 8 0 0 4
157 488
218 488
218 611
231 611
6 1 18 0 0 4224 0 12 9 0 0 4
157 479
225 479
225 537
233 537
5 1 19 0 0 4224 0 12 6 0 0 2
157 470
233 470
2 1 20 0 0 4224 0 6 18 0 0 4
269 470
271 470
271 470
269 470
4 1 21 0 0 4224 0 14 11 0 0 3
335 129
453 129
453 67
5 1 22 0 0 8320 0 17 10 0 0 3
335 369
503 369
503 66
5 2 23 0 0 8320 0 16 10 0 0 3
335 282
497 282
497 66
5 3 24 0 0 4224 0 15 10 0 0 3
335 195
491 195
491 66
5 4 25 0 0 4224 0 14 10 0 0 3
335 111
485 111
485 66
1 3 8 0 0 128 0 4 17 0 0 4
43 432
241 432
241 387
269 387
4 3 26 0 0 12416 0 15 14 0 0 5
335 213
353 213
353 156
269 156
269 129
4 3 27 0 0 12416 0 16 15 0 0 5
335 300
353 300
353 242
269 242
269 213
4 3 28 0 0 12416 0 17 16 0 0 5
335 387
353 387
353 329
269 329
269 300
1 1 29 0 0 4224 0 13 17 0 0 3
127 70
127 369
269 369
2 1 30 0 0 4224 0 13 16 0 0 3
121 70
121 282
269 282
3 1 31 0 0 8320 0 13 15 0 0 3
115 70
115 195
269 195
4 1 32 0 0 8320 0 13 14 0 0 3
109 70
109 111
269 111
4 8 16 0 0 0 0 12 12 0 0 6
87 497
83 497
83 512
165 512
165 497
157 497
1 3 33 0 0 4224 0 5 12 0 0 2
40 488
87 488
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
