CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
370 80 3 160 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
10
12 Hex Display~
7 595 66 0 16 19
10 2 3 4 5 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
5130 0 0
2
5.89855e-315 0
0
12 Hex Display~
7 421 71 0 16 19
10 6 7 8 9 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
391 0 0
2
5.89855e-315 0
0
5 4071~
219 518 204 0 3 22
0 11 12 10
0
0 0 624 180
4 4071
-7 -24 21 -16
3 U4A
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
3124 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 508 146 0 3 22
0 13 14 11
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U3D
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
3421 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 586 145 0 3 22
0 5 5 14
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U3C
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
8157 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 427 207 0 3 22
0 7 7 13
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U3B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
5572 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 586 207 0 3 22
0 5 3 12
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U3A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
8901 0 0
2
5.89855e-315 0
0
7 Pulser~
4 505 359 0 10 12
0 16 17 15 18 0 0 5 5 6
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7361 0 0
2
5.89855e-315 0
0
6 74LS93
109 585 275 0 8 17
0 10 10 15 2 5 4 3 2
0
0 0 4848 0
6 74LS93
-21 -35 21 -27
2 U2
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
4747 0 0
2
5.89855e-315 0
0
6 74LS93
109 424 275 0 8 17
0 11 11 5 6 9 8 7 6
0
0 0 4848 0
6 74LS93
-21 -35 21 -27
2 U1
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
972 0 0
2
5.89855e-315 0
0
26
8 1 2 0 0 8320 0 9 1 0 0 5
617 293
661 293
661 113
604 113
604 90
7 2 3 0 0 8320 0 9 1 0 0 5
617 284
656 284
656 108
598 108
598 90
6 3 4 0 0 8320 0 9 1 0 0 5
617 275
651 275
651 103
592 103
592 90
5 4 5 0 0 8192 0 9 1 0 0 5
617 266
646 266
646 98
586 98
586 90
8 1 6 0 0 8320 0 10 2 0 0 5
456 293
475 293
475 118
430 118
430 95
7 2 7 0 0 8320 0 10 2 0 0 5
456 284
475 284
475 113
424 113
424 95
6 3 8 0 0 8320 0 10 2 0 0 5
456 275
475 275
475 108
418 108
418 95
5 4 9 0 0 8320 0 10 2 0 0 5
456 266
470 266
470 103
412 103
412 95
0 2 10 0 0 8192 0 0 9 10 0 3
517 266
517 275
553 275
3 1 10 0 0 4224 0 3 9 0 0 3
491 204
491 266
553 266
3 1 11 0 0 8192 0 4 3 0 0 6
481 146
479 146
479 231
556 231
556 213
537 213
2 3 12 0 0 4224 0 3 7 0 0 6
537 195
610 195
610 227
556 227
556 207
559 207
3 2 11 0 0 8320 0 4 10 0 0 4
481 146
373 146
373 275
392 275
3 1 11 0 0 0 0 4 10 0 0 4
481 146
378 146
378 266
392 266
3 1 13 0 0 12416 0 6 4 0 0 6
400 207
398 207
398 126
541 126
541 155
526 155
3 2 14 0 0 4224 0 5 4 0 0 4
559 145
536 145
536 137
526 137
5 2 5 0 0 0 0 9 5 0 0 4
617 266
641 266
641 136
604 136
5 1 5 0 0 0 0 9 5 0 0 4
617 266
636 266
636 154
604 154
7 2 7 0 0 0 0 10 6 0 0 4
456 284
465 284
465 198
445 198
7 1 7 0 0 0 0 10 6 0 0 4
456 284
460 284
460 216
445 216
7 2 3 0 0 0 0 9 7 0 0 4
617 284
631 284
631 198
604 198
5 1 5 0 0 0 0 9 7 0 0 4
617 266
621 266
621 216
604 216
8 4 6 0 0 0 0 10 10 0 0 6
456 293
460 293
460 308
373 308
373 293
386 293
5 3 5 0 0 12416 0 9 10 0 0 6
617 266
626 266
626 313
378 313
378 284
386 284
8 4 2 0 0 0 0 9 9 0 0 6
617 293
621 293
621 308
534 308
534 293
547 293
3 3 15 0 0 8320 0 8 9 0 0 4
529 350
539 350
539 284
547 284
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
426 389 599 413
432 394 592 410
20 DIVIDE BY 27 COUNTER
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
