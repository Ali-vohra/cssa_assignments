CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
70 30 30 120 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
14
13 Logic Switch~
5 313 61 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8157 0 0
2
43332 0
0
13 Logic Switch~
5 129 307 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5572 0 0
2
43332 0
0
13 Logic Switch~
5 130 267 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8901 0 0
2
43332 0
0
13 Logic Switch~
5 131 172 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7361 0 0
2
43332 0
0
13 Logic Switch~
5 131 133 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4747 0 0
2
43332 0
0
9 2-In AND~
219 252 264 0 3 22
0 8 7 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
972 0 0
2
43332 0
0
9 2-In AND~
219 252 214 0 3 22
0 11 7 10
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3472 0 0
2
43332 0
0
6 74LS83
105 457 230 0 14 29
0 3 3 6 12 3 3 3 10 3
14 4 5 9 15
0
0 0 4848 0
5 74F83
-18 -60 17 -52
2 U2
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 0 0 0 0
1 U
9998 0 0
2
43332 0
0
9 2-In AND~
219 252 166 0 3 22
0 8 13 12
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3536 0 0
2
43332 0
0
14 Logic Display~
6 960 189 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4597 0 0
2
43332 0
0
14 Logic Display~
6 961 262 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3835 0 0
2
43332 0
0
14 Logic Display~
6 965 343 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3670 0 0
2
43332 0
0
14 Logic Display~
6 963 419 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5616 0 0
2
43332 0
0
9 2-In AND~
219 252 113 0 3 22
0 11 13 2
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
9323 0 0
2
43332 0
0
21
3 1 2 0 0 4224 0 14 13 0 0 5
273 113
933 113
933 448
963 448
963 437
1 5 3 0 0 8192 0 1 8 0 0 4
325 61
387 61
387 230
425 230
1 1 3 0 0 0 0 1 8 0 0 4
325 61
402 61
402 194
425 194
11 1 4 0 0 4224 0 8 10 0 0 3
489 230
960 230
960 207
1 2 3 0 0 0 0 1 8 0 0 4
325 61
412 61
412 203
425 203
1 6 3 0 0 8192 0 1 8 0 0 4
325 61
392 61
392 239
425 239
12 1 5 0 0 4224 0 8 11 0 0 5
489 239
943 239
943 288
961 288
961 280
1 7 3 0 0 8192 0 1 8 0 0 4
325 61
397 61
397 248
425 248
3 3 6 0 0 4224 0 6 8 0 0 4
273 264
402 264
402 212
425 212
1 2 7 0 0 4096 0 3 6 0 0 4
142 267
205 267
205 273
228 273
1 1 8 0 0 8320 0 5 6 0 0 4
143 133
205 133
205 255
228 255
13 1 9 0 0 4224 0 8 12 0 0 5
489 248
949 248
949 369
965 369
965 361
1 9 3 0 0 8320 0 1 8 0 0 4
325 61
407 61
407 275
425 275
3 8 10 0 0 4224 0 7 8 0 0 4
273 214
412 214
412 257
425 257
1 2 7 0 0 4224 0 3 7 0 0 4
142 267
210 267
210 223
228 223
1 1 11 0 0 4096 0 4 7 0 0 4
143 172
210 172
210 205
228 205
3 4 12 0 0 4224 0 9 8 0 0 4
273 166
417 166
417 221
425 221
1 2 13 0 0 8192 0 2 9 0 0 4
141 307
220 307
220 175
228 175
1 1 8 0 0 0 0 5 9 0 0 4
143 133
210 133
210 157
228 157
1 2 13 0 0 8320 0 2 14 0 0 4
141 307
215 307
215 122
228 122
1 1 11 0 0 4224 0 4 14 0 0 4
143 172
220 172
220 104
228 104
9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
478 429 623 450
486 436 614 451
16 2 BIT MULTIPLIER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
968 178 1003 199
977 185 993 200
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
966 252 1001 273
975 259 991 274
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
970 333 1003 354
978 340 994 355
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
969 409 1002 430
977 416 993 431
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
74 287 111 311
84 295 100 311
2 B0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
77 247 114 271
87 255 103 271
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
77 157 114 181
87 165 103 181
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
77 113 114 137
87 121 103 137
2 A1
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
