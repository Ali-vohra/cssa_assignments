CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
21
13 Logic Switch~
5 561 251 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43354 0
0
13 Logic Switch~
5 30 384 0 1 11
0 24
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
43354 0
0
13 Logic Switch~
5 31 432 0 1 11
0 25
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89861e-315 0
0
13 Logic Switch~
5 28 488 0 1 11
0 26
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
5.89861e-315 0
0
12 Hex Display~
7 195 330 0 18 19
10 2 3 4 5 0 0 0 0 0
0 1 0 1 1 1 1 1 6
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
8157 0 0
2
43354 0
0
8 2-In OR~
219 757 159 0 3 22
0 8 7 6
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U12A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
5572 0 0
2
43354 0
0
12 Hex Display~
7 850 42 0 18 19
10 9 10 11 12 0 0 0 0 0
0 1 0 1 1 0 1 1 5
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
8901 0 0
2
43354 0
0
12 Hex Display~
7 805 43 0 18 19
10 6 58 59 60 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 0 0 0 0
4 DISP
7361 0 0
2
43354 0
0
8 3-In OR~
219 519 182 0 4 22
0 23 7 22 14
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U7A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 2 0
1 U
4747 0 0
2
43354 0
0
9 2-In AND~
219 412 235 0 3 22
0 21 19 22
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
972 0 0
2
43354 0
0
9 2-In AND~
219 413 143 0 3 22
0 21 20 23
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3472 0 0
2
43354 0
0
6 74LS90
107 125 470 0 10 21
0 24 24 25 25 26 2 5 4 3
2
0
0 0 4848 0
6 74LS90
-21 -51 21 -43
2 U5
-7 -52 7 -44
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 0 0 0 0
1 U
9998 0 0
2
43354 0
0
8 Hex Key~
166 118 46 0 11 12
0 30 31 32 33 0 0 0 0 0
9 57
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3536 0 0
2
5.89861e-315 0
0
2 FA
94 302 111 0 5 11
0 33 5 27 7 21
2 FA
1 0 688 0
0
2 U1
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 1 0 0 0
1 U
4597 0 0
2
5.89859e-315 0
0
2 FA
94 302 195 0 5 11
0 32 4 28 27 20
2 FA
2 0 688 0
0
2 U2
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 1 0 0 0
1 U
3835 0 0
2
5.89859e-315 0
0
2 FA
94 302 282 0 5 11
0 31 3 29 28 19
2 FA
3 0 688 0
0
2 U3
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 1 0 0 0
1 U
3670 0 0
2
5.89859e-315 0
0
2 FA
94 302 369 0 5 11
0 30 2 24 29 18
2 FA
4 0 688 0
0
2 U4
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 1 0 0 0
1 U
5616 0 0
2
5.89859e-315 0
0
2 FA
94 662 111 0 5 11
0 21 13 15 8 12
2 FA
5 0 688 0
0
2 U8
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
9323 0 0
2
43334.9 0
0
2 FA
94 661 192 0 5 11
0 20 14 16 15 11
2 FA
6 0 688 0
0
2 U9
-7 -29 7 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
317 0 0
2
43334.9 0
0
2 FA
94 660 282 0 5 11
0 19 14 17 16 10
2 FA
7 0 688 0
0
3 U10
-11 -29 10 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
3108 0 0
2
43334.9 0
0
2 FA
94 659 369 0 5 11
0 18 13 13 17 9
2 FA
8 0 688 0
0
3 U11
-11 -29 10 -21
0
0
0
0
0
0
11

0 1 2 3 4 6 1 2 3 4
6 0
0 0 0 0 0 0 0 0
1 U
4299 0 0
2
43334.9 0
0
48
10 1 2 0 0 8320 0 12 5 0 0 3
157 497
204 497
204 354
9 2 3 0 0 8192 0 12 5 0 0 3
157 479
198 479
198 354
8 3 4 0 0 8192 0 12 5 0 0 3
157 461
192 461
192 354
7 4 5 0 0 8192 0 12 5 0 0 3
157 443
186 443
186 354
3 1 6 0 0 8320 0 6 8 0 0 3
790 159
814 159
814 67
4 2 7 0 0 12416 0 14 6 0 0 8
335 129
370 129
370 207
624 207
624 229
736 229
736 168
744 168
4 1 8 0 0 4224 0 18 6 0 0 4
695 129
736 129
736 150
744 150
5 1 9 0 0 8320 0 21 7 0 0 3
692 369
859 369
859 66
5 2 10 0 0 8320 0 20 7 0 0 3
693 282
853 282
853 66
5 3 11 0 0 4224 0 19 7 0 0 3
694 192
847 192
847 66
5 4 12 0 0 4224 0 18 7 0 0 3
695 111
841 111
841 66
1 3 13 0 0 8320 0 1 21 0 0 4
573 251
603 251
603 387
626 387
1 2 13 0 0 0 0 1 21 0 0 4
573 251
613 251
613 378
626 378
1 2 13 0 0 0 0 1 18 0 0 4
573 251
606 251
606 120
629 120
4 2 14 0 0 8320 0 9 20 0 0 4
552 182
609 182
609 291
627 291
4 2 14 0 0 0 0 9 19 0 0 4
552 182
615 182
615 201
628 201
4 3 15 0 0 12416 0 19 18 0 0 6
694 210
699 210
699 143
621 143
621 129
629 129
4 3 16 0 0 12416 0 20 19 0 0 6
693 300
698 300
698 224
620 224
620 210
628 210
4 3 17 0 0 12416 0 21 20 0 0 6
692 387
697 387
697 314
619 314
619 300
627 300
5 1 18 0 0 4224 0 17 21 0 0 2
335 369
626 369
5 1 19 0 0 4224 0 16 20 0 0 2
335 282
627 282
5 1 20 0 0 4224 0 15 19 0 0 6
335 195
502 195
502 202
620 202
620 192
628 192
5 1 21 0 0 4224 0 14 18 0 0 2
335 111
629 111
4 2 7 0 0 128 0 14 9 0 0 4
335 129
385 129
385 182
507 182
3 3 22 0 0 4224 0 10 9 0 0 4
433 235
498 235
498 191
506 191
3 1 23 0 0 4224 0 11 9 0 0 4
434 143
498 143
498 173
506 173
5 2 19 0 0 0 0 16 10 0 0 4
335 282
380 282
380 244
388 244
5 1 21 0 0 0 0 14 10 0 0 4
335 111
375 111
375 226
388 226
5 2 20 0 0 0 0 15 11 0 0 4
335 195
381 195
381 152
389 152
5 1 21 0 0 0 0 14 11 0 0 4
335 111
381 111
381 134
389 134
1 3 24 0 0 4224 0 2 17 0 0 4
42 384
241 384
241 387
269 387
10 2 2 0 0 128 0 12 17 0 0 4
157 497
246 497
246 378
269 378
9 2 3 0 0 8320 0 12 16 0 0 4
157 479
251 479
251 291
269 291
8 2 4 0 0 8320 0 12 15 0 0 4
157 461
256 461
256 204
269 204
7 2 5 0 0 8320 0 12 14 0 0 4
157 443
261 443
261 120
269 120
1 2 24 0 0 0 0 2 12 0 0 4
42 384
64 384
64 452
93 452
1 1 24 0 0 0 0 2 12 0 0 4
42 384
69 384
69 443
93 443
1 3 25 0 0 4096 0 3 12 0 0 4
43 432
74 432
74 461
93 461
1 4 25 0 0 8320 0 3 12 0 0 4
43 432
79 432
79 470
93 470
10 6 2 0 0 0 0 12 12 0 0 6
157 497
161 497
161 512
79 512
79 497
87 497
1 5 26 0 0 4224 0 4 12 0 0 2
40 488
87 488
4 3 27 0 0 12416 0 15 14 0 0 5
335 213
353 213
353 156
269 156
269 129
4 3 28 0 0 12416 0 16 15 0 0 5
335 300
353 300
353 242
269 242
269 213
4 3 29 0 0 12416 0 17 16 0 0 5
335 387
353 387
353 329
269 329
269 300
1 1 30 0 0 4224 0 13 17 0 0 3
127 70
127 369
269 369
2 1 31 0 0 4224 0 13 16 0 0 3
121 70
121 282
269 282
3 1 32 0 0 8320 0 13 15 0 0 3
115 70
115 195
269 195
4 1 33 0 0 8320 0 13 14 0 0 3
109 70
109 111
269 111
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
