CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
240 40 7 140 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
15
12 Hex Display~
7 756 85 0 18 19
10 2 3 4 5 0 0 0 0 0
0 1 0 1 1 1 1 1 6
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
5130 0 0
2
5.89855e-315 0
0
12 Hex Display~
7 528 91 0 18 19
10 6 7 8 9 0 0 0 0 0
0 1 1 0 1 1 0 1 2
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
391 0 0
2
5.89855e-315 0
0
12 Hex Display~
7 296 96 0 16 19
10 10 11 12 13 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3124 0 0
2
5.89855e-315 0
0
5 4071~
219 665 252 0 3 22
0 15 16 14
0
0 0 608 180
4 4071
-7 -24 21 -16
3 U7B
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 4 0
1 U
3421 0 0
2
5.89855e-315 0
0
5 4071~
219 427 254 0 3 22
0 18 15 17
0
0 0 608 180
4 4071
-7 -24 21 -16
3 U7A
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
8157 0 0
2
5.89855e-315 0
0
5 4073~
219 293 188 0 4 22
0 21 20 19 15
0
0 0 608 180
4 4073
-7 -24 21 -16
3 U6A
-13 -25 8 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 3 0
1 U
5572 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 757 192 0 3 22
0 5 2 19
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U5A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
8901 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 523 197 0 3 22
0 7 6 20
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U4D
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
7361 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 294 256 0 3 22
0 11 11 21
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U4C
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
4747 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 522 256 0 3 22
0 9 7 18
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U4B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
972 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 757 254 0 3 22
0 5 3 16
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U4A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3472 0 0
2
5.89855e-315 0
0
7 Pulser~
4 672 415 0 10 12
0 23 24 22 25 0 0 5 5 1
8
0
0 0 4640 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
9998 0 0
2
5.89855e-315 0
0
6 74LS93
109 756 318 0 8 17
0 14 14 22 2 5 4 3 2
0
0 0 4832 0
6 74LS93
-21 -35 21 -27
2 U3
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
3536 0 0
2
5.89855e-315 0
0
6 74LS93
109 521 321 0 8 17
0 17 17 5 6 9 8 7 6
0
0 0 4832 0
6 74LS93
-21 -35 21 -27
2 U2
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
4597 0 0
2
5.89855e-315 0
0
6 74LS93
109 293 322 0 8 17
0 15 15 9 10 13 12 11 10
0
0 0 4832 0
6 74LS93
-21 -35 21 -27
2 U1
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
3835 0 0
2
5.89855e-315 0
0
41
8 1 2 0 0 8320 0 13 1 0 0 5
788 336
832 336
832 132
765 132
765 109
7 2 3 0 0 8320 0 13 1 0 0 5
788 327
827 327
827 127
759 127
759 109
6 3 4 0 0 8320 0 13 1 0 0 5
788 318
822 318
822 122
753 122
753 109
5 4 5 0 0 8192 0 13 1 0 0 5
788 309
817 309
817 117
747 117
747 109
8 1 6 0 0 8320 0 14 2 0 0 5
553 339
597 339
597 138
537 138
537 115
7 2 7 0 0 8320 0 14 2 0 0 5
553 330
592 330
592 133
531 133
531 115
6 3 8 0 0 8320 0 14 2 0 0 5
553 321
587 321
587 128
525 128
525 115
5 4 9 0 0 8192 0 14 2 0 0 5
553 312
582 312
582 123
519 123
519 115
8 1 10 0 0 8320 0 15 3 0 0 5
325 340
354 340
354 143
305 143
305 120
7 2 11 0 0 8320 0 15 3 0 0 5
325 331
349 331
349 138
299 138
299 120
6 3 12 0 0 8320 0 15 3 0 0 5
325 322
344 322
344 133
293 133
293 120
5 4 13 0 0 8320 0 15 3 0 0 5
325 313
339 313
339 128
287 128
287 120
3 2 14 0 0 8320 0 4 13 0 0 3
638 252
638 318
724 318
3 1 14 0 0 0 0 4 13 0 0 3
638 252
638 309
724 309
4 1 15 0 0 12416 0 6 4 0 0 6
266 188
255 188
255 281
706 281
706 261
684 261
2 3 16 0 0 4224 0 4 11 0 0 4
684 243
724 243
724 254
730 254
0 2 17 0 0 8192 0 0 14 18 0 3
423 312
423 321
489 321
3 1 17 0 0 8320 0 5 14 0 0 3
400 254
400 312
489 312
3 1 18 0 0 12416 0 10 5 0 0 4
495 256
473 256
473 263
446 263
4 2 15 0 0 0 0 6 5 0 0 6
266 188
260 188
260 276
468 276
468 245
446 245
4 2 15 0 0 0 0 6 15 0 0 4
266 188
242 188
242 322
261 322
4 1 15 0 0 0 0 6 15 0 0 4
266 188
247 188
247 313
261 313
3 3 19 0 0 12416 0 7 6 0 0 4
730 192
547 192
547 179
311 179
3 2 20 0 0 4224 0 8 6 0 0 4
496 197
326 197
326 188
311 188
3 1 21 0 0 8320 0 9 6 0 0 6
267 256
264 256
264 168
321 168
321 197
311 197
8 2 2 0 0 0 0 13 7 0 0 4
788 336
812 336
812 183
775 183
5 1 5 0 0 0 0 13 7 0 0 4
788 309
807 309
807 201
775 201
8 2 6 0 0 0 0 14 8 0 0 4
553 339
577 339
577 188
541 188
7 1 7 0 0 0 0 14 8 0 0 4
553 330
572 330
572 206
541 206
7 2 11 0 0 0 0 15 9 0 0 4
325 331
334 331
334 247
312 247
7 1 11 0 0 0 0 15 9 0 0 4
325 331
329 331
329 265
312 265
7 2 7 0 0 0 0 14 10 0 0 4
553 330
567 330
567 247
540 247
5 1 9 0 0 0 0 14 10 0 0 4
553 312
557 312
557 265
540 265
7 2 3 0 0 0 0 13 11 0 0 4
788 327
802 327
802 245
775 245
5 1 5 0 0 0 0 13 11 0 0 4
788 309
792 309
792 263
775 263
8 4 10 0 0 0 0 15 15 0 0 6
325 340
329 340
329 355
242 355
242 340
255 340
5 3 9 0 0 12416 0 14 15 0 0 6
553 312
562 312
562 364
247 364
247 331
255 331
8 4 6 0 0 0 0 14 14 0 0 6
553 339
557 339
557 359
470 359
470 339
483 339
5 3 5 0 0 12416 0 13 14 0 0 6
788 309
797 309
797 354
475 354
475 330
483 330
8 4 2 0 0 0 0 13 13 0 0 6
788 336
792 336
792 351
705 351
705 336
718 336
3 3 22 0 0 8320 0 12 13 0 0 4
696 406
710 406
710 327
718 327
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
472 449 655 473
479 454 647 470
21 3 BIT COUNTER IC 7493
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
