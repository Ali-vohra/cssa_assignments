CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
220 50 30 170 10
176 80 1534 843
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
17
13 Logic Switch~
5 617 212 0 1 11
0 6
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9323 0 0
2
43319.7 0
0
13 Logic Switch~
5 369 291 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
317 0 0
2
43319.7 0
0
14 Logic Display~
6 924 282 0 1 2
10 30
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 0 0 0 0
1 L
3108 0 0
2
43319.7 0
0
12 Hex Display~
7 916 164 0 16 19
10 2 3 4 5 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
4299 0 0
2
43319.7 0
0
5 4049~
219 497 341 0 2 22
0 8 7
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 3 0
1 U
9672 0 0
2
43319.7 0
0
5 4030~
219 590 466 0 3 22
0 13 7 9
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U4D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 2 0
1 U
7876 0 0
2
43319.7 0
0
5 4030~
219 592 413 0 3 22
0 14 7 10
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U4C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
6369 0 0
2
43319.7 0
0
5 4030~
219 591 362 0 3 22
0 15 7 11
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U4B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
9172 0 0
2
43319.7 0
0
5 4030~
219 591 312 0 3 22
0 16 7 12
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U4A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
7100 0 0
2
43319.7 0
0
6 74LS83
105 738 252 0 14 29
0 6 6 6 6 12 11 10 9 7
5 4 3 2 31
0
0 0 4848 0
5 74F83
-18 -60 17 -52
2 U3
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 0 0 0 0
1 U
3820 0 0
2
43319.7 0
0
9 Inverter~
13 296 415 0 2 22
0 22 18
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
7678 0 0
2
43319.7 3
0
9 Inverter~
13 295 382 0 2 22
0 23 19
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
961 0 0
2
43319.7 4
0
9 Inverter~
13 294 350 0 2 22
0 24 20
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
3178 0 0
2
43319.7 5
0
9 Inverter~
13 293 318 0 2 22
0 25 21
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3409 0 0
2
43319.7 6
0
8 Hex Key~
166 245 141 0 11 12
0 22 23 24 25 0 0 0 0 0
0 48
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3951 0 0
2
43319.7 7
0
8 Hex Key~
166 337 143 0 11 12
0 26 27 28 29 0 0 0 0 0
0 48
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
8885 0 0
2
43319.7 8
0
6 74LS83
105 477 257 0 14 29
0 29 28 27 26 21 20 19 18 17
16 15 14 13 8
0
0 0 4848 0
5 74F83
-18 -60 17 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
3780 0 0
2
43319.7 9
0
36
14 1 0 0 0 0 0 10 3 0 0 5
770 297
912 297
912 308
924 308
924 300
13 1 2 0 0 4224 0 10 4 0 0 5
770 270
902 270
902 196
925 196
925 188
12 2 3 0 0 4224 0 10 4 0 0 3
770 261
919 261
919 188
11 3 4 0 0 4224 0 10 4 0 0 3
770 252
913 252
913 188
10 4 5 0 0 4224 0 10 4 0 0 3
770 243
907 243
907 188
1 4 6 0 0 4096 0 1 10 0 0 4
629 212
683 212
683 243
706 243
1 3 6 0 0 4096 0 1 10 0 0 4
629 212
688 212
688 234
706 234
1 2 6 0 0 4096 0 1 10 0 0 4
629 212
693 212
693 225
706 225
1 1 6 0 0 4224 0 1 10 0 0 4
629 212
698 212
698 216
706 216
2 9 7 0 0 4224 0 5 10 0 0 4
518 341
678 341
678 297
706 297
2 2 7 0 0 0 0 5 6 0 0 4
518 341
536 341
536 475
574 475
2 2 7 0 0 0 0 5 7 0 0 4
518 341
543 341
543 422
576 422
2 2 7 0 0 0 0 5 8 0 0 4
518 341
547 341
547 371
575 371
2 2 7 0 0 0 0 5 9 0 0 4
518 341
567 341
567 321
575 321
14 1 8 0 0 8320 0 17 5 0 0 6
509 302
522 302
522 356
474 356
474 341
482 341
3 8 9 0 0 8320 0 6 10 0 0 4
623 466
683 466
683 279
706 279
3 7 10 0 0 8320 0 7 10 0 0 4
625 413
688 413
688 270
706 270
3 6 11 0 0 8320 0 8 10 0 0 4
624 362
693 362
693 261
706 261
3 5 12 0 0 4224 0 9 10 0 0 4
624 312
698 312
698 252
706 252
13 1 13 0 0 8320 0 17 6 0 0 4
509 275
551 275
551 457
574 457
12 1 14 0 0 8320 0 17 7 0 0 4
509 266
558 266
558 404
576 404
11 1 15 0 0 8320 0 17 8 0 0 4
509 257
562 257
562 353
575 353
10 1 16 0 0 4224 0 17 9 0 0 4
509 248
567 248
567 303
575 303
1 9 17 0 0 4224 0 2 17 0 0 4
381 291
417 291
417 302
445 302
2 8 18 0 0 8320 0 11 17 0 0 4
317 415
422 415
422 284
445 284
2 7 19 0 0 4224 0 12 17 0 0 4
316 382
427 382
427 275
445 275
2 6 20 0 0 4224 0 13 17 0 0 4
315 350
432 350
432 266
445 266
2 5 21 0 0 4224 0 14 17 0 0 4
314 318
437 318
437 257
445 257
1 1 22 0 0 4224 0 15 11 0 0 3
254 165
254 415
281 415
2 1 23 0 0 4224 0 15 12 0 0 3
248 165
248 382
280 382
3 1 24 0 0 4224 0 15 13 0 0 3
242 165
242 350
279 350
4 1 25 0 0 4224 0 15 14 0 0 3
236 165
236 318
278 318
1 4 26 0 0 8320 0 16 17 0 0 3
346 167
346 248
445 248
2 3 27 0 0 8320 0 16 17 0 0 3
340 167
340 239
445 239
3 2 28 0 0 8320 0 16 17 0 0 3
334 167
334 230
445 230
4 1 29 0 0 8320 0 16 17 0 0 3
328 167
328 221
445 221
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
395 59 592 83
405 67 581 83
22 BINARY SUBTRACTOR(2'S)
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
