CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
40 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
24
13 Logic Switch~
5 152 429 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43331.5 0
0
13 Logic Switch~
5 151 214 0 10 11
0 27 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
391 0 0
2
43331.5 0
0
9 2-In AND~
219 1006 146 0 3 22
0 4 3 2
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
3124 0 0
2
43331.5 0
0
9 Inverter~
13 933 361 0 2 22
0 6 3
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 5 0
1 U
3421 0 0
2
43331.5 0
0
9 Inverter~
13 926 207 0 2 22
0 5 4
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 5 0
1 U
8157 0 0
2
43331.5 0
0
5 4073~
219 808 231 0 4 22
0 10 7 8 5
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 4 0
1 U
5572 0 0
2
43331.5 0
0
9 Inverter~
13 707 494 0 2 22
0 9 8
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
8901 0 0
2
43331.5 0
0
9 Inverter~
13 577 400 0 2 22
0 11 10
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
7361 0 0
2
43331.5 0
0
9 2-In AND~
219 675 274 0 3 22
0 13 12 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
4747 0 0
2
43331.5 0
0
14 Logic Display~
6 1122 143 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
972 0 0
2
43331.5 0
0
14 Logic Display~
6 1123 252 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3472 0 0
2
43331.5 0
0
14 Logic Display~
6 1123 353 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9998 0 0
2
43331.5 0
0
8 2-In OR~
219 871 388 0 3 22
0 9 11 6
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3536 0 0
2
43331.5 0
0
8 2-In OR~
219 670 428 0 3 22
0 14 15 9
0
0 0 624 270
6 74LS32
-21 -24 21 -16
3 U5A
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
4597 0 0
2
43331.5 0
0
9 2-In AND~
219 709 365 0 3 22
0 16 13 14
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U4B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3835 0 0
2
43331.5 0
0
9 2-In AND~
219 639 366 0 3 22
0 17 13 15
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U4A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3670 0 0
2
43331.5 0
0
6 74LS83
105 518 323 0 14 29
0 26 25 24 23 22 21 20 19 18
13 17 16 12 11
0
0 0 4848 0
5 74F83
-18 -60 17 -52
2 U3
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 0 0 0 0
1 U
5616 0 0
2
43331.5 0
0
8 Hex Key~
166 330 78 0 11 12
0 23 24 25 26 0 0 0 0 0
4 52
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
9323 0 0
2
43331.5 0
0
6 74LS83
105 329 325 0 14 29
0 27 18 27 18 31 30 29 28 18
22 21 20 19 36
0
0 0 4848 0
5 74F83
-18 -60 17 -52
2 U2
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 0 0 0 0
1 U
317 0 0
2
43331.5 0
0
9 Inverter~
13 148 388 0 2 22
0 32 28
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
3108 0 0
2
43331.5 0
0
9 Inverter~
13 149 348 0 2 22
0 33 29
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
4299 0 0
2
43331.5 0
0
9 Inverter~
13 149 309 0 2 22
0 34 30
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
9672 0 0
2
43331.5 0
0
9 Inverter~
13 149 271 0 2 22
0 35 31
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
7876 0 0
2
43331.5 0
0
8 Hex Key~
166 61 79 0 11 12
0 32 33 34 35 0 0 0 0 0
5 53
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
6369 0 0
2
43331.5 0
0
44
3 1 2 0 0 4224 0 3 10 0 0 5
1027 146
1110 146
1110 169
1122 169
1122 161
2 2 3 0 0 8320 0 4 3 0 0 4
954 361
969 361
969 155
982 155
2 1 4 0 0 8320 0 5 3 0 0 4
947 207
974 207
974 137
982 137
4 1 5 0 0 4096 0 6 5 0 0 4
829 231
903 231
903 207
911 207
3 1 6 0 0 8192 0 13 4 0 0 4
904 388
910 388
910 361
918 361
4 1 5 0 0 4224 0 6 11 0 0 5
829 231
1110 231
1110 278
1123 278
1123 270
3 2 7 0 0 4224 0 9 6 0 0 4
696 274
776 274
776 231
784 231
2 3 8 0 0 8320 0 7 6 0 0 5
728 494
748 494
748 299
784 299
784 240
3 1 9 0 0 4096 0 14 7 0 0 3
673 458
673 494
692 494
2 1 10 0 0 4224 0 8 6 0 0 5
598 400
598 236
696 236
696 222
784 222
14 1 11 0 0 8192 0 17 8 0 0 4
550 368
554 368
554 400
562 400
13 2 12 0 0 4224 0 17 9 0 0 4
550 341
618 341
618 283
651 283
10 1 13 0 0 4096 0 17 9 0 0 4
550 314
643 314
643 265
651 265
3 1 6 0 0 4224 0 13 12 0 0 3
904 388
1123 388
1123 371
14 2 11 0 0 12416 0 17 13 0 0 5
550 368
612 368
612 468
858 468
858 397
3 1 9 0 0 8320 0 14 13 0 0 5
673 458
673 455
850 455
850 379
858 379
3 1 14 0 0 8320 0 15 14 0 0 4
707 388
707 397
682 397
682 412
3 2 15 0 0 8320 0 16 14 0 0 4
637 389
637 397
664 397
664 412
12 1 16 0 0 4224 0 17 15 0 0 3
550 332
716 332
716 343
10 2 13 0 0 4224 0 17 15 0 0 3
550 314
698 314
698 343
11 1 17 0 0 4224 0 17 16 0 0 3
550 323
646 323
646 344
10 2 13 0 0 0 0 17 16 0 0 3
550 314
628 314
628 344
1 9 18 0 0 4224 0 1 17 0 0 4
164 429
478 429
478 368
486 368
13 8 19 0 0 4224 0 19 17 0 0 4
361 343
478 343
478 350
486 350
12 7 20 0 0 4224 0 19 17 0 0 4
361 334
478 334
478 341
486 341
11 6 21 0 0 4224 0 19 17 0 0 4
361 325
478 325
478 332
486 332
10 5 22 0 0 4224 0 19 17 0 0 4
361 316
478 316
478 323
486 323
1 4 23 0 0 4224 0 18 17 0 0 5
339 102
339 255
463 255
463 314
486 314
2 3 24 0 0 4224 0 18 17 0 0 5
333 102
333 260
468 260
468 305
486 305
3 2 25 0 0 4224 0 18 17 0 0 5
327 102
327 265
473 265
473 296
486 296
4 1 26 0 0 4224 0 18 17 0 0 5
321 102
321 270
478 270
478 287
486 287
1 4 18 0 0 0 0 1 19 0 0 4
164 429
269 429
269 316
297 316
1 2 18 0 0 0 0 1 19 0 0 4
164 429
274 429
274 298
297 298
1 9 18 0 0 0 0 1 19 0 0 4
164 429
289 429
289 370
297 370
1 3 27 0 0 4096 0 2 19 0 0 4
163 214
279 214
279 307
297 307
1 1 27 0 0 4224 0 2 19 0 0 4
163 214
284 214
284 289
297 289
2 8 28 0 0 4224 0 20 19 0 0 4
169 388
283 388
283 352
297 352
2 7 29 0 0 4224 0 21 19 0 0 4
170 348
279 348
279 343
297 343
2 6 30 0 0 4224 0 22 19 0 0 4
170 309
283 309
283 334
297 334
2 5 31 0 0 4224 0 23 19 0 0 4
170 271
289 271
289 325
297 325
1 1 32 0 0 4224 0 24 20 0 0 3
70 103
70 388
133 388
2 1 33 0 0 4224 0 24 21 0 0 3
64 103
64 348
134 348
3 1 34 0 0 4224 0 24 22 0 0 3
58 103
58 309
134 309
4 1 35 0 0 4224 0 24 23 0 0 3
52 103
52 271
134 271
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
487 543 668 567
497 551 657 567
20 BCD COMPARATOR (9'S)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
47 12 76 36
57 20 65 36
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
317 13 346 37
327 21 335 37
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1127 129 1172 153
1137 137 1161 153
3 A<B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1129 235 1174 259
1139 243 1163 259
3 A=B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1129 341 1174 365
1139 349 1163 365
3 A>B
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
