CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
220 50 30 140 10
176 80 1534 843
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
23
13 Logic Switch~
5 617 212 0 1 11
0 16
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89857e-315 0
0
13 Logic Switch~
5 369 291 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.89857e-315 0
0
9 2-In AND~
219 759 420 0 3 22
0 4 3 2
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3124 0 0
2
43319.7 0
0
9 Inverter~
13 707 527 0 2 22
0 4 5
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
3421 0 0
2
43319.7 0
0
8 4-In OR~
219 594 532 0 5 22
0 9 8 7 6 4
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U6A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 4 0
1 U
8157 0 0
2
43319.7 0
0
14 Logic Display~
6 932 535 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5572 0 0
2
43319.7 0
0
14 Logic Display~
6 931 465 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8901 0 0
2
43319.7 0
0
14 Logic Display~
6 928 394 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7361 0 0
2
43319.7 0
0
14 Logic Display~
6 924 282 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4747 0 0
2
5.89857e-315 0
0
12 Hex Display~
7 916 164 0 18 19
10 12 13 14 15 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
972 0 0
2
5.89857e-315 0
0
5 4049~
219 497 341 0 2 22
0 3 10
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 3 0
1 U
3472 0 0
2
5.89857e-315 0
0
5 4030~
219 590 466 0 3 22
0 6 10 17
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U4D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 2 0
1 U
9998 0 0
2
5.89857e-315 0
0
5 4030~
219 592 413 0 3 22
0 7 10 18
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U4C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
3536 0 0
2
5.89857e-315 0
0
5 4030~
219 591 362 0 3 22
0 8 10 19
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U4B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
4597 0 0
2
5.89857e-315 0
0
5 4030~
219 591 312 0 3 22
0 9 10 20
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U4A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
3835 0 0
2
5.89857e-315 0
0
6 74LS83
105 738 252 0 14 29
0 16 16 16 16 20 19 18 17 10
15 14 13 12 11
0
0 0 4848 0
5 74F83
-18 -60 17 -52
2 U3
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
3670 0 0
2
5.89857e-315 0
0
9 Inverter~
13 296 415 0 2 22
0 26 22
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
5616 0 0
2
5.89857e-315 5.32571e-315
0
9 Inverter~
13 295 382 0 2 22
0 27 23
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
9323 0 0
2
5.89857e-315 5.34643e-315
0
9 Inverter~
13 294 350 0 2 22
0 28 24
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
317 0 0
2
5.89857e-315 5.3568e-315
0
9 Inverter~
13 293 318 0 2 22
0 29 25
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3108 0 0
2
5.89857e-315 5.36716e-315
0
8 Hex Key~
166 245 141 0 11 12
0 26 27 28 29 0 0 0 0 0
3 51
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
4299 0 0
2
5.89857e-315 5.37752e-315
0
8 Hex Key~
166 337 143 0 11 12
0 30 31 32 33 0 0 0 0 0
2 50
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
9672 0 0
2
5.89857e-315 5.38788e-315
0
6 74LS83
105 477 257 0 14 29
0 33 32 31 30 25 24 23 22 21
9 8 7 6 3
0
0 0 4848 0
5 74F83
-18 -60 17 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
7876 0 0
2
5.89857e-315 5.39306e-315
0
46
3 1 2 0 0 4224 0 3 8 0 0 3
780 420
928 420
928 412
14 2 3 0 0 12416 0 23 3 0 0 6
509 302
572 302
572 433
727 433
727 429
735 429
5 1 4 0 0 8320 0 5 3 0 0 4
627 532
678 532
678 411
735 411
2 1 5 0 0 4224 0 4 7 0 0 5
728 527
920 527
920 491
931 491
931 483
5 1 4 0 0 0 0 5 4 0 0 4
627 532
684 532
684 527
692 527
13 4 6 0 0 8320 0 23 5 0 0 4
509 275
524 275
524 546
577 546
12 3 7 0 0 8320 0 23 5 0 0 4
509 266
539 266
539 537
577 537
2 11 8 0 0 8320 0 5 23 0 0 4
577 528
528 528
528 257
509 257
10 1 9 0 0 8320 0 23 5 0 0 4
509 248
554 248
554 519
577 519
2 1 10 0 0 4224 0 11 6 0 0 5
518 341
944 341
944 561
932 561
932 553
14 1 11 0 0 4224 0 16 9 0 0 5
770 297
912 297
912 308
924 308
924 300
13 1 12 0 0 4224 0 16 10 0 0 5
770 270
902 270
902 196
925 196
925 188
12 2 13 0 0 4224 0 16 10 0 0 3
770 261
919 261
919 188
11 3 14 0 0 4224 0 16 10 0 0 3
770 252
913 252
913 188
10 4 15 0 0 4224 0 16 10 0 0 3
770 243
907 243
907 188
1 4 16 0 0 4096 0 1 16 0 0 4
629 212
683 212
683 243
706 243
1 3 16 0 0 4096 0 1 16 0 0 4
629 212
688 212
688 234
706 234
1 2 16 0 0 4096 0 1 16 0 0 4
629 212
693 212
693 225
706 225
1 1 16 0 0 4224 0 1 16 0 0 4
629 212
698 212
698 216
706 216
2 9 10 0 0 128 0 11 16 0 0 4
518 341
678 341
678 297
706 297
2 2 10 0 0 0 0 11 12 0 0 4
518 341
536 341
536 475
574 475
2 2 10 0 0 0 0 11 13 0 0 4
518 341
543 341
543 422
576 422
2 2 10 0 0 0 0 11 14 0 0 4
518 341
547 341
547 371
575 371
2 2 10 0 0 0 0 11 15 0 0 4
518 341
567 341
567 321
575 321
14 1 3 0 0 128 0 23 11 0 0 6
509 302
522 302
522 356
474 356
474 341
482 341
3 8 17 0 0 8320 0 12 16 0 0 4
623 466
683 466
683 279
706 279
3 7 18 0 0 8320 0 13 16 0 0 4
625 413
688 413
688 270
706 270
3 6 19 0 0 8320 0 14 16 0 0 4
624 362
693 362
693 261
706 261
3 5 20 0 0 4224 0 15 16 0 0 4
624 312
698 312
698 252
706 252
13 1 6 0 0 128 0 23 12 0 0 4
509 275
551 275
551 457
574 457
12 1 7 0 0 128 0 23 13 0 0 4
509 266
558 266
558 404
576 404
11 1 8 0 0 128 0 23 14 0 0 4
509 257
562 257
562 353
575 353
10 1 9 0 0 128 0 23 15 0 0 4
509 248
567 248
567 303
575 303
1 9 21 0 0 4224 0 2 23 0 0 4
381 291
417 291
417 302
445 302
2 8 22 0 0 8320 0 17 23 0 0 4
317 415
422 415
422 284
445 284
2 7 23 0 0 4224 0 18 23 0 0 4
316 382
427 382
427 275
445 275
2 6 24 0 0 4224 0 19 23 0 0 4
315 350
432 350
432 266
445 266
2 5 25 0 0 4224 0 20 23 0 0 4
314 318
437 318
437 257
445 257
1 1 26 0 0 4224 0 21 17 0 0 3
254 165
254 415
281 415
2 1 27 0 0 4224 0 21 18 0 0 3
248 165
248 382
280 382
3 1 28 0 0 4224 0 21 19 0 0 3
242 165
242 350
279 350
4 1 29 0 0 4224 0 21 20 0 0 3
236 165
236 318
278 318
1 4 30 0 0 8320 0 22 23 0 0 3
346 167
346 248
445 248
2 3 31 0 0 8320 0 22 23 0 0 3
340 167
340 239
445 239
3 2 32 0 0 8320 0 22 23 0 0 3
334 167
334 230
445 230
4 1 33 0 0 8320 0 22 23 0 0 3
328 167
328 221
445 221
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
947 524 984 548
953 529 977 545
3 A<B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
947 456 984 480
953 461 977 477
3 A=B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
947 383 984 407
953 388 977 404
3 A>B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
395 59 592 83
405 67 581 83
22 BINARY SUBTRACTOR(2'S)
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
