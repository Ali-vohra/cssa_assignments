CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
250 60 5 160 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
8
13 Logic Switch~
5 444 219 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43329.9 0
0
9 2-In AND~
219 543 164 0 3 22
0 5 6 4
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U3B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
391 0 0
2
43329.9 0
0
9 2-In AND~
219 306 169 0 3 22
0 4 7 3
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U3A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3124 0 0
2
43329.9 0
0
12 Hex Display~
7 677 105 0 18 19
10 5 11 6 12 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3421 0 0
2
43329.9 0
0
12 Hex Display~
7 406 112 0 18 19
10 8 9 7 10 0 0 0 0 0
0 1 1 0 1 1 0 1 2
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
8157 0 0
2
43329.9 0
0
7 Pulser~
4 426 351 0 10 12
0 14 15 13 16 0 0 5 5 3
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
5572 0 0
2
43329.9 0
0
6 74LS90
107 540 250 0 10 21
0 2 2 3 3 13 5 12 6 11
5
0
0 0 4848 0
6 74LS90
-21 -51 21 -43
2 U2
-7 -52 7 -44
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 0 0 0 0
1 U
8901 0 0
2
43329.9 0
0
6 74LS93
109 307 263 0 8 17
0 3 3 12 8 10 7 9 8
0
0 0 4848 0
6 74LS93
-21 -35 21 -27
2 U1
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 0 0 0 0
1 U
7361 0 0
2
43329.9 0
0
22
1 2 2 0 0 4096 0 1 7 0 0 4
456 219
489 219
489 232
508 232
1 1 2 0 0 4224 0 1 7 0 0 4
456 219
494 219
494 223
508 223
3 4 3 0 0 12416 0 3 7 0 0 6
279 169
250 169
250 311
479 311
479 250
508 250
3 3 3 0 0 0 0 3 7 0 0 6
279 169
265 169
265 306
484 306
484 241
508 241
3 2 3 0 0 0 0 3 8 0 0 4
279 169
256 169
256 263
275 263
3 1 3 0 0 0 0 3 8 0 0 4
279 169
261 169
261 254
275 254
3 1 4 0 0 4224 0 2 3 0 0 4
516 164
334 164
334 178
324 178
10 1 5 0 0 8192 0 7 2 0 0 4
572 277
591 277
591 173
561 173
2 8 6 0 0 8192 0 2 7 0 0 4
561 155
585 155
585 241
572 241
6 2 7 0 0 8192 0 8 3 0 0 4
339 263
343 263
343 160
324 160
8 1 8 0 0 8320 0 8 5 0 0 3
339 281
415 281
415 136
7 2 9 0 0 8320 0 8 5 0 0 3
339 272
409 272
409 136
6 3 7 0 0 8320 0 8 5 0 0 3
339 263
403 263
403 136
5 4 10 0 0 8320 0 8 5 0 0 3
339 254
397 254
397 136
10 1 5 0 0 8320 0 7 4 0 0 3
572 277
686 277
686 129
9 2 11 0 0 8320 0 7 4 0 0 3
572 259
680 259
680 129
8 3 6 0 0 8320 0 7 4 0 0 3
572 241
674 241
674 129
7 4 12 0 0 4096 0 7 4 0 0 3
572 223
668 223
668 129
8 4 8 0 0 0 0 8 8 0 0 6
339 281
343 281
343 301
256 301
256 281
269 281
7 3 12 0 0 12416 0 7 8 0 0 6
572 223
581 223
581 296
261 296
261 272
269 272
10 6 5 0 0 0 0 7 7 0 0 6
572 277
576 277
576 292
489 292
489 277
502 277
3 5 13 0 0 8320 0 6 7 0 0 4
450 342
494 342
494 268
502 268
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
337 405 520 429
344 410 512 426
21 45 COUNTER (COMBINED)
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
