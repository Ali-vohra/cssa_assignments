CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 50 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
80
13 Logic Switch~
5 60 401 0 10 11
0 71 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 60 351 0 10 11
0 69 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 60 302 0 10 11
0 67 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 60 254 0 10 11
0 65 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 57 167 0 10 11
0 70 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 57 121 0 10 11
0 68 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 57 73 0 10 11
0 66 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 58 32 0 10 11
0 64 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7361 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 1304 667 0 3 22
0 4 5 3
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U13D
-15 -4 13 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 16 0
1 U
4747 0 0
2
43337.5 0
0
9 2-In XOR~
219 1296 617 0 3 22
0 4 5 2
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U12D
-3 -4 25 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 15 0
1 U
972 0 0
2
43337.5 0
0
9 2-In AND~
219 1305 562 0 3 22
0 7 8 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U13C
-16 -4 12 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 16 0
1 U
3472 0 0
2
43337.5 0
0
9 2-In XOR~
219 1298 510 0 3 22
0 7 8 4
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U12C
-3 -5 25 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 15 0
1 U
9998 0 0
2
43337.5 0
0
9 2-In AND~
219 1105 877 0 3 22
0 12 13 10
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U13B
-16 -4 12 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 16 0
1 U
3536 0 0
2
43337.5 0
0
9 2-In XOR~
219 1098 827 0 3 22
0 13 12 9
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U12B
-3 -4 25 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 15 0
1 U
4597 0 0
2
43337.5 0
0
9 2-In AND~
219 1107 773 0 3 22
0 14 15 11
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U13A
-16 -3 12 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 16 0
1 U
3835 0 0
2
43337.5 0
0
9 2-In XOR~
219 1099 723 0 3 22
0 14 15 12
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U12A
-3 -4 25 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 15 0
1 U
3670 0 0
2
43337.5 0
0
9 2-In AND~
219 1109 666 0 3 22
0 17 18 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U11D
-16 -3 12 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 14 0
1 U
5616 0 0
2
43337.5 0
0
9 2-In XOR~
219 1101 617 0 3 22
0 18 17 13
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U10D
-3 -4 25 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 13 0
1 U
9323 0 0
2
43337.5 0
0
9 2-In AND~
219 1110 563 0 3 22
0 20 21 19
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U11C
-16 -3 12 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 14 0
1 U
317 0 0
2
43337.5 0
0
9 2-In XOR~
219 1102 513 0 3 22
0 20 21 18
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U10C
-3 -3 25 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 13 0
1 U
3108 0 0
2
43337.5 0
0
9 2-In AND~
219 862 993 0 3 22
0 23 24 17
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U11B
-16 -4 12 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 14 0
1 U
4299 0 0
2
43337.5 0
0
9 2-In XOR~
219 854 939 0 3 22
0 23 24 22
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U10B
-3 -4 25 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 13 0
1 U
9672 0 0
2
43337.5 0
0
9 2-In AND~
219 865 884 0 3 22
0 27 28 25
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U11A
-16 -3 12 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 14 0
1 U
7876 0 0
2
43337.5 0
0
9 2-In XOR~
219 859 836 0 3 22
0 27 28 24
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U10A
-3 -4 25 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 13 0
1 U
6369 0 0
2
43337.5 0
0
9 2-In AND~
219 869 778 0 3 22
0 29 30 26
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9D
-12 -4 9 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 12 0
1 U
9172 0 0
2
43337.5 0
0
9 2-In XOR~
219 862 727 0 3 22
0 29 30 28
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6D
0 -4 21 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 11 0
1 U
7100 0 0
2
43337.5 0
0
9 2-In AND~
219 872 672 0 3 22
0 32 33 31
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9C
-13 -4 8 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 12 0
1 U
3820 0 0
2
43337.5 0
0
9 2-In XOR~
219 864 623 0 3 22
0 32 33 23
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6C
0 -3 21 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
7678 0 0
2
43337.5 0
0
9 2-In AND~
219 873 568 0 3 22
0 35 36 34
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9B
-12 -3 9 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 12 0
1 U
961 0 0
2
43337.5 0
0
9 2-In XOR~
219 868 515 0 3 22
0 35 36 33
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6B
0 -4 21 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
3178 0 0
2
43337.5 0
0
9 2-In AND~
219 582 1001 0 3 22
0 39 38 32
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9A
-13 -3 8 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 12 0
1 U
3409 0 0
2
43337.5 0
0
9 2-In XOR~
219 574 946 0 3 22
0 38 39 37
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U6A
0 -4 21 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
3951 0 0
2
43337.5 0
0
9 2-In AND~
219 583 885 0 3 22
0 41 42 40
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5D
-12 -4 9 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 10 0
1 U
8885 0 0
2
43337.5 0
0
9 2-In XOR~
219 577 832 0 3 22
0 42 41 39
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U4D
0 -3 21 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 9 0
1 U
3780 0 0
2
43337.5 0
0
9 2-In AND~
219 586 774 0 3 22
0 44 45 43
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5C
-13 -3 8 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 10 0
1 U
9265 0 0
2
43337.5 0
0
9 2-In XOR~
219 578 724 0 3 22
0 45 44 41
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U4C
0 -4 21 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
9442 0 0
2
43337.5 0
0
9 2-In AND~
219 587 671 0 3 22
0 47 48 46
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5B
-13 -4 8 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 10 0
1 U
9424 0 0
2
43337.5 0
0
9 2-In XOR~
219 580 624 0 3 22
0 47 48 38
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U4B
-1 -4 20 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
9968 0 0
2
43337.5 0
0
9 2-In AND~
219 588 573 0 3 22
0 50 51 49
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -3 9 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
9281 0 0
2
43337.5 0
0
9 2-In XOR~
219 581 524 0 3 22
0 50 51 47
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U4A
0 -4 21 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
8464 0 0
2
43337.5 0
0
9 2-In AND~
219 319 793 0 3 22
0 54 53 51
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U27D
-16 -3 12 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 8 0
1 U
7168 0 0
2
43337.5 0
0
9 2-In XOR~
219 313 739 0 3 22
0 54 53 52
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U2D
0 -3 21 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
3171 0 0
2
43337.5 0
0
9 2-In AND~
219 321 683 0 3 22
0 57 58 55
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U27C
-16 -3 12 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 8 0
1 U
4139 0 0
2
43337.5 0
0
9 2-In XOR~
219 313 634 0 3 22
0 57 58 54
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U2C
0 -3 21 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
6435 0 0
2
43337.5 0
0
9 2-In AND~
219 322 580 0 3 22
0 59 60 56
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U27B
-16 -4 12 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
5283 0 0
2
43337.5 0
0
9 2-In XOR~
219 315 532 0 3 22
0 59 60 58
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U2B
0 -3 21 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
6874 0 0
2
43337.5 0
0
9 2-In AND~
219 181 579 0 3 22
0 61 62 53
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U27A
-15 -4 13 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
5305 0 0
2
43337.5 0
0
9 2-In XOR~
219 175 532 0 3 22
0 62 61 72
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U2A
0 -4 21 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
34 0 0
2
43337.5 0
0
14 Logic Display~
6 1490 1114 0 1 2
10 63
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
969 0 0
2
5.89859e-315 0
0
14 Logic Display~
6 1384 1116 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8402 0 0
2
5.89859e-315 0
0
14 Logic Display~
6 1173 1117 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3751 0 0
2
5.89859e-315 0
0
14 Logic Display~
6 944 1120 0 1 2
10 22
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4292 0 0
2
5.89859e-315 0
0
14 Logic Display~
6 687 1120 0 1 2
10 37
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6118 0 0
2
5.89859e-315 0
0
14 Logic Display~
6 418 1118 0 1 2
10 52
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
34 0 0
2
5.89859e-315 0
0
14 Logic Display~
6 287 1121 0 1 2
10 72
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6357 0 0
2
5.89859e-315 0
0
14 Logic Display~
6 149 1122 0 1 2
10 73
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
319 0 0
2
5.89859e-315 0
0
8 2-In OR~
219 1406 545 0 3 22
0 6 3 63
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U20D
-4 -4 24 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
3976 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 1302 444 0 3 22
0 64 65 5
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U14D
-14 -10 14 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
7634 0 0
2
5.89859e-315 0
0
8 2-In OR~
219 1196 714 0 3 22
0 11 10 7
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U20C
-4 -4 24 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
523 0 0
2
5.89859e-315 0
0
8 2-In OR~
219 1196 552 0 3 22
0 19 16 8
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U20B
-4 -4 24 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
6748 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 1125 445 0 3 22
0 65 66 14
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U14C
-15 -11 13 -3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
6901 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 1083 446 0 3 22
0 67 64 15
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U14B
-15 -10 13 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
842 0 0
2
5.89859e-315 0
0
8 2-In OR~
219 968 716 0 3 22
0 26 25 20
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U20A
-3 -4 25 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
3277 0 0
2
5.89859e-315 0
0
8 2-In OR~
219 970 558 0 3 22
0 34 31 21
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7D
-1 -4 20 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
4212 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 907 445 0 3 22
0 65 68 27
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U14A
-15 -10 13 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
4720 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 866 446 0 3 22
0 67 66 30
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U8D
-12 -10 9 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
5551 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 826 446 0 3 22
0 69 64 29
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U8C
-12 -9 9 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
6986 0 0
2
5.89859e-315 0
0
8 2-In OR~
219 703 713 0 3 22
0 43 40 36
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7C
0 -2 21 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
8745 0 0
2
5.89859e-315 0
0
8 2-In OR~
219 705 561 0 3 22
0 49 46 35
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7B
-1 -4 20 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
9592 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 654 447 0 3 22
0 65 70 42
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U8B
-12 -9 9 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
8748 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 614 447 0 3 22
0 67 68 44
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U8A
-12 -9 9 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
7168 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 572 448 0 3 22
0 69 66 45
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3D
-11 -9 10 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
631 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 530 449 0 3 22
0 71 64 48
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3C
-11 -8 10 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
9466 0 0
2
5.89859e-315 0
0
8 2-In OR~
219 426 644 0 3 22
0 56 55 50
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U7A
-1 -3 20 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3266 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 366 450 0 3 22
0 67 70 57
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3B
-12 -9 9 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
7693 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 320 451 0 3 22
0 69 68 60
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U3A
-12 -9 9 -1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3723 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 275 451 0 3 22
0 71 66 59
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1D
-12 -8 9 0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
3440 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 207 450 0 3 22
0 69 70 61
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1C
-12 -6 9 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
6263 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 158 451 0 3 22
0 71 68 62
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1B
-12 -6 9 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
4900 0 0
2
5.89859e-315 0
0
9 2-In AND~
219 108 450 0 3 22
0 71 70 73
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U1A
-12 -5 9 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
8783 0 0
2
5.89859e-315 0
0
144
3 1 2 0 0 8320 0 10 50 0 0 5
1329 617
1349 617
1349 1159
1384 1159
1384 1134
3 2 3 0 0 8320 0 9 57 0 0 4
1325 667
1380 667
1380 554
1393 554
0 1 4 0 0 4096 0 0 9 5 0 3
1253 608
1253 658
1280 658
0 2 5 0 0 4096 0 0 9 6 0 3
1246 626
1246 676
1280 676
3 1 4 0 0 12416 0 12 10 0 0 6
1331 510
1341 510
1341 590
1253 590
1253 608
1280 608
3 2 5 0 0 8320 0 58 10 0 0 4
1300 467
1233 467
1233 626
1280 626
3 1 6 0 0 4224 0 11 57 0 0 4
1326 562
1385 562
1385 536
1393 536
0 1 7 0 0 4096 0 0 11 10 0 3
1258 501
1258 553
1281 553
0 2 8 0 0 4096 0 0 11 11 0 3
1247 519
1247 571
1281 571
3 1 7 0 0 8320 0 59 12 0 0 4
1229 714
1238 714
1238 501
1282 501
3 2 8 0 0 8320 0 60 12 0 0 3
1229 552
1229 519
1282 519
3 1 9 0 0 8320 0 14 51 0 0 5
1131 827
1141 827
1141 1159
1173 1159
1173 1135
3 2 10 0 0 8320 0 13 59 0 0 4
1126 877
1170 877
1170 723
1183 723
3 1 11 0 0 8320 0 15 59 0 0 4
1128 773
1175 773
1175 705
1183 705
0 1 12 0 0 8192 0 0 13 18 0 3
1042 836
1042 868
1081 868
0 2 13 0 0 4096 0 0 13 17 0 3
1033 818
1033 886
1081 886
3 1 13 0 0 8320 0 18 14 0 0 6
1134 617
1146 617
1146 805
1033 805
1033 818
1082 818
3 2 12 0 0 12416 0 16 14 0 0 6
1132 723
1151 723
1151 798
1042 798
1042 836
1082 836
0 1 14 0 0 4096 0 0 15 21 0 3
1054 714
1054 764
1083 764
0 2 15 0 0 4096 0 0 15 22 0 3
1042 732
1042 782
1083 782
3 1 14 0 0 8320 0 61 16 0 0 6
1123 468
1156 468
1156 695
1054 695
1054 714
1083 714
3 2 15 0 0 8320 0 62 16 0 0 4
1081 469
1042 469
1042 732
1083 732
3 2 16 0 0 8320 0 17 60 0 0 4
1130 666
1175 666
1175 561
1183 561
0 1 17 0 0 8192 0 0 17 27 0 3
1028 626
1028 657
1085 657
0 2 18 0 0 4096 0 0 17 26 0 3
1021 608
1021 675
1085 675
3 1 18 0 0 12416 0 20 18 0 0 6
1135 513
1146 513
1146 590
1021 590
1021 608
1085 608
3 2 17 0 0 8320 0 21 18 0 0 4
883 993
1007 993
1007 626
1085 626
3 1 19 0 0 4224 0 19 60 0 0 4
1131 563
1170 563
1170 543
1183 543
0 1 20 0 0 4096 0 0 19 31 0 3
1067 504
1067 554
1086 554
0 2 21 0 0 4096 0 0 19 32 0 3
1054 522
1054 572
1086 572
3 1 20 0 0 8320 0 63 20 0 0 4
1001 716
1013 716
1013 504
1086 504
3 2 21 0 0 8320 0 64 20 0 0 3
1003 558
1003 522
1086 522
3 1 22 0 0 8320 0 22 52 0 0 5
887 939
893 939
893 1159
944 1159
944 1138
0 1 23 0 0 4096 0 0 21 36 0 3
793 930
793 984
838 984
0 2 24 0 0 4096 0 0 21 37 0 3
802 948
802 1002
838 1002
3 1 23 0 0 8320 0 28 22 0 0 6
897 623
913 623
913 918
793 918
793 930
838 930
3 2 24 0 0 12416 0 24 22 0 0 6
892 836
917 836
917 912
802 912
802 948
838 948
3 2 25 0 0 8320 0 23 63 0 0 4
886 884
942 884
942 725
955 725
3 1 26 0 0 8320 0 25 63 0 0 4
890 778
947 778
947 707
955 707
0 1 27 0 0 4096 0 0 23 42 0 3
794 826
794 875
841 875
0 2 28 0 0 8192 0 0 23 43 0 3
787 845
787 893
841 893
3 1 27 0 0 4224 0 65 24 0 0 5
905 468
905 813
794 813
794 827
843 827
3 2 28 0 0 12416 0 26 24 0 0 6
895 727
928 727
928 804
787 804
787 845
843 845
0 1 29 0 0 8192 0 0 25 47 0 3
773 718
773 769
845 769
0 2 30 0 0 8192 0 0 25 46 0 3
767 735
767 787
845 787
3 2 30 0 0 12416 0 66 26 0 0 5
864 469
864 478
767 478
767 736
846 736
3 1 29 0 0 8320 0 67 26 0 0 4
824 469
773 469
773 718
846 718
3 2 31 0 0 8320 0 27 64 0 0 4
893 672
949 672
949 567
957 567
0 1 32 0 0 4096 0 0 27 51 0 3
813 614
813 663
848 663
0 2 33 0 0 4096 0 0 27 52 0 3
802 632
802 681
848 681
3 1 32 0 0 8320 0 31 28 0 0 4
603 1001
780 1001
780 614
848 614
3 2 33 0 0 12416 0 30 28 0 0 6
901 515
921 515
921 597
802 597
802 632
848 632
3 1 34 0 0 4224 0 29 64 0 0 4
894 568
944 568
944 549
957 549
0 1 35 0 0 4096 0 0 29 57 0 3
831 506
831 559
849 559
0 2 36 0 0 4096 0 0 29 56 0 3
810 524
810 577
849 577
3 2 36 0 0 8320 0 68 30 0 0 4
736 713
787 713
787 524
852 524
3 1 35 0 0 12416 0 69 30 0 0 4
738 561
793 561
793 506
852 506
3 1 37 0 0 8320 0 32 53 0 0 5
607 946
651 946
651 1159
687 1159
687 1138
0 2 38 0 0 4096 0 0 31 61 0 3
492 937
492 1010
558 1010
0 1 39 0 0 8192 0 0 31 62 0 3
498 953
498 992
558 992
3 1 38 0 0 8320 0 38 32 0 0 6
613 624
644 624
644 921
492 921
492 937
558 937
3 2 39 0 0 12416 0 34 32 0 0 6
610 832
638 832
638 914
498 914
498 955
558 955
3 2 40 0 0 8320 0 33 68 0 0 4
604 885
677 885
677 722
690 722
0 1 41 0 0 8192 0 0 33 67 0 3
507 841
507 876
559 876
0 2 42 0 0 4096 0 0 33 66 0 3
498 823
498 894
559 894
3 1 42 0 0 4224 0 70 34 0 0 5
652 470
652 812
498 812
498 823
561 823
3 2 41 0 0 12416 0 36 34 0 0 6
611 724
638 724
638 803
507 803
507 841
561 841
3 1 43 0 0 4224 0 35 68 0 0 4
607 774
682 774
682 704
690 704
0 1 44 0 0 8192 0 0 35 71 0 3
461 733
461 765
562 765
0 2 45 0 0 8192 0 0 35 72 0 3
483 714
483 783
562 783
3 2 44 0 0 12416 0 71 36 0 0 5
612 470
612 491
461 491
461 733
562 733
3 1 45 0 0 12416 0 72 36 0 0 5
570 471
570 481
483 481
483 715
562 715
3 2 46 0 0 8320 0 37 69 0 0 4
608 671
684 671
684 570
692 570
0 1 47 0 0 4096 0 0 37 76 0 3
516 615
516 662
563 662
0 2 48 0 0 8192 0 0 37 77 0 3
507 633
507 680
563 680
3 1 47 0 0 12416 0 40 38 0 0 6
614 524
638 524
638 600
516 600
516 615
564 615
3 2 48 0 0 8320 0 73 38 0 0 4
528 472
507 472
507 633
564 633
3 1 49 0 0 4224 0 39 69 0 0 4
609 573
679 573
679 552
692 552
0 1 50 0 0 4096 0 0 39 82 0 3
533 515
533 564
564 564
0 2 51 0 0 4096 0 0 39 81 0 3
517 533
517 582
564 582
3 2 51 0 0 8320 0 41 40 0 0 4
340 793
494 793
494 533
565 533
3 1 50 0 0 8320 0 74 40 0 0 4
459 644
472 644
472 515
565 515
3 1 52 0 0 8320 0 42 54 0 0 5
346 739
372 739
372 1158
418 1158
418 1136
0 2 53 0 0 4096 0 0 41 87 0 3
255 748
255 802
295 802
0 1 54 0 0 4096 0 0 41 86 0 3
278 730
278 784
295 784
3 1 54 0 0 12416 0 44 42 0 0 6
346 634
372 634
372 712
278 712
278 730
297 730
3 2 53 0 0 8320 0 47 42 0 0 4
202 579
221 579
221 748
297 748
3 2 55 0 0 4224 0 43 74 0 0 4
342 683
405 683
405 653
413 653
3 1 56 0 0 4224 0 45 74 0 0 4
343 580
405 580
405 635
413 635
0 1 57 0 0 4096 0 0 43 92 0 3
265 625
265 674
297 674
0 2 58 0 0 4096 0 0 43 93 0 3
258 643
258 692
297 692
3 1 57 0 0 4224 0 75 44 0 0 5
364 473
364 604
265 604
265 625
297 625
3 2 58 0 0 12416 0 46 44 0 0 6
348 532
380 532
380 609
258 609
258 643
297 643
0 1 59 0 0 4096 0 0 45 96 0 3
273 523
273 571
298 571
0 2 60 0 0 4096 0 0 45 97 0 3
258 540
258 589
298 589
3 1 59 0 0 4224 0 77 46 0 0 3
273 474
273 523
299 523
3 2 60 0 0 8320 0 76 46 0 0 5
318 474
318 500
258 500
258 541
299 541
0 1 61 0 0 4096 0 0 47 101 0 3
141 541
141 570
157 570
0 2 62 0 0 4224 0 0 47 100 0 3
132 523
132 588
157 588
3 1 62 0 0 0 0 79 48 0 0 5
156 474
156 491
132 491
132 523
159 523
3 2 61 0 0 8320 0 78 48 0 0 5
205 473
205 502
141 502
141 541
159 541
3 1 63 0 0 8320 0 57 49 0 0 5
1439 545
1465 545
1465 1159
1490 1159
1490 1132
1 0 64 0 0 4096 0 58 0 0 144 2
1309 422
1309 32
2 0 65 0 0 4096 0 58 0 0 140 2
1291 422
1291 254
1 0 65 0 0 4096 0 61 0 0 140 2
1132 423
1132 254
2 0 66 0 0 4096 0 61 0 0 143 2
1114 423
1114 73
1 0 67 0 0 4096 0 62 0 0 139 2
1090 424
1090 302
2 0 64 0 0 4096 0 62 0 0 144 2
1072 424
1072 32
1 0 65 0 0 0 0 65 0 0 140 2
914 423
914 254
2 0 68 0 0 4096 0 65 0 0 142 2
896 423
896 121
1 0 67 0 0 0 0 66 0 0 139 2
873 424
873 302
2 0 66 0 0 4096 0 66 0 0 143 2
855 424
855 73
1 0 69 0 0 4096 0 67 0 0 138 2
833 424
833 351
2 0 64 0 0 0 0 67 0 0 144 2
815 424
815 32
1 0 65 0 0 4096 0 70 0 0 140 2
661 425
661 254
2 0 70 0 0 4096 0 70 0 0 141 2
643 425
643 167
1 0 67 0 0 4096 0 71 0 0 139 2
621 425
621 302
2 0 68 0 0 4096 0 71 0 0 142 2
603 425
603 121
1 0 69 0 0 4096 0 72 0 0 138 2
579 426
579 351
2 0 66 0 0 4096 0 72 0 0 143 2
561 426
561 73
1 0 71 0 0 4096 0 73 0 0 137 2
537 427
537 401
2 0 64 0 0 4096 0 73 0 0 144 2
519 427
519 32
1 0 67 0 0 4096 0 75 0 0 139 2
373 428
373 302
2 0 70 0 0 4096 0 75 0 0 141 2
355 428
355 167
1 0 69 0 0 4096 0 76 0 0 138 2
327 429
327 351
2 0 68 0 0 4096 0 76 0 0 142 2
309 429
309 121
1 0 71 0 0 4096 0 77 0 0 137 2
282 429
282 401
2 0 66 0 0 4096 0 77 0 0 143 2
264 429
264 73
3 1 72 0 0 8320 0 48 55 0 0 5
208 532
229 532
229 1158
287 1158
287 1139
1 0 69 0 0 0 0 78 0 0 138 2
214 428
214 351
2 0 70 0 0 0 0 78 0 0 141 2
196 428
196 167
1 0 71 0 0 0 0 79 0 0 137 2
165 429
165 401
2 0 68 0 0 0 0 79 0 0 142 2
147 429
147 121
3 1 73 0 0 4224 0 80 56 0 0 4
106 473
106 1158
149 1158
149 1140
2 0 70 0 0 0 0 80 0 0 141 2
97 428
97 167
1 0 71 0 0 0 0 80 0 0 137 2
115 428
115 401
1 0 71 0 0 4224 0 1 0 0 0 2
72 401
1552 401
1 0 69 0 0 4224 0 2 0 0 0 2
72 351
1552 351
1 0 67 0 0 4224 0 3 0 0 0 2
72 302
1551 302
1 0 65 0 0 4224 0 4 0 0 0 2
72 254
1551 254
1 0 70 0 0 4224 0 5 0 0 0 2
69 167
1551 167
1 0 68 0 0 4224 0 6 0 0 0 2
69 121
1551 121
1 0 66 0 0 4224 0 7 0 0 0 2
69 73
1552 73
1 0 64 0 0 4224 0 8 0 0 0 2
70 32
1552 32
16
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
7 10 44 34
17 18 33 34
2 A3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
7 51 44 75
17 59 33 75
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
8 99 45 123
18 107 34 123
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
8 144 45 168
18 152 34 168
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
11 230 48 254
21 238 37 254
2 B3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
12 283 49 307
22 291 38 307
2 B2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
10 332 47 356
20 340 36 356
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
10 377 47 401
20 385 36 401
2 B0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
127 1057 170 1072
141 1069 155 1080
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
262 1060 307 1075
277 1071 291 1082
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
395 1060 440 1075
410 1071 424 1082
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
665 1063 708 1078
679 1075 693 1086
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
922 1064 965 1079
936 1075 950 1086
2 S4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1150 1062 1195 1077
1165 1074 1179 1085
2 S5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1361 1061 1406 1076
1376 1072 1390 1083
2 S6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1469 1061 1514 1076
1484 1072 1498 1083
2 S7
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
