CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1534 843
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
22
13 Logic Switch~
5 121 353 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3409 0 0
2
43318.7 0
0
13 Logic Switch~
5 123 302 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3951 0 0
2
43318.7 0
0
13 Logic Switch~
5 119 206 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8885 0 0
2
43318.7 0
0
13 Logic Switch~
5 120 156 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3780 0 0
2
43318.7 0
0
14 Logic Display~
6 911 322 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9265 0 0
2
43318.7 0
0
14 Logic Display~
6 911 222 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9442 0 0
2
43318.7 0
0
14 Logic Display~
6 908 121 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9424 0 0
2
43318.7 0
0
5 4071~
219 730 342 0 3 22
0 5 6 2
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U4B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 4 0
1 U
9968 0 0
2
43318.7 0
0
9 2-In AND~
219 586 351 0 3 22
0 8 7 6
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
9281 0 0
2
43318.7 0
0
9 2-In AND~
219 366 360 0 3 22
0 10 9 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
8464 0 0
2
43318.7 0
0
9 2-In AND~
219 364 305 0 3 22
0 12 11 5
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
7168 0 0
2
43318.7 0
0
9 2-In AND~
219 739 246 0 3 22
0 8 13 3
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
3171 0 0
2
43318.7 0
0
10 2-In XNOR~
219 440 290 0 3 22
0 14 9 13
0
0 0 624 0
4 4077
-7 -24 21 -16
3 U3B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 3 0
1 U
4139 0 0
2
43318.7 0
0
5 4071~
219 730 156 0 3 22
0 16 15 4
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
6435 0 0
2
43318.7 0
0
9 2-In AND~
219 598 162 0 3 22
0 8 17 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
5283 0 0
2
43318.7 0
0
10 2-In XNOR~
219 441 163 0 3 22
0 18 11 8
0
0 0 624 0
4 4077
-7 -24 21 -16
3 U3A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
6874 0 0
2
43318.7 0
0
9 2-In AND~
219 353 200 0 3 22
0 14 19 17
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
5305 0 0
2
43318.7 0
0
9 2-In AND~
219 354 146 0 3 22
0 18 20 15
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
34 0 0
2
43318.7 0
0
9 Inverter~
13 233 350 0 2 22
0 9 19
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
969 0 0
2
43318.7 0
0
9 Inverter~
13 233 294 0 2 22
0 14 10
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
8402 0 0
2
43318.7 0
0
9 Inverter~
13 234 198 0 2 22
0 11 20
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
3751 0 0
2
43318.7 0
0
9 Inverter~
13 232 153 0 2 22
0 18 12
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
4292 0 0
2
43318.7 0
0
29
3 1 2 0 0 4224 0 8 5 0 0 5
763 342
899 342
899 348
911 348
911 340
3 1 3 0 0 4224 0 12 6 0 0 3
760 246
911 246
911 240
3 1 4 0 0 4224 0 14 7 0 0 3
763 156
908 156
908 139
3 1 5 0 0 12416 0 11 8 0 0 6
385 305
420 305
420 371
709 371
709 333
717 333
3 2 6 0 0 4224 0 9 8 0 0 2
607 351
717 351
3 2 7 0 0 4224 0 10 9 0 0 2
387 360
562 360
3 1 8 0 0 8320 0 16 9 0 0 6
480 163
492 163
492 326
435 326
435 342
562 342
1 2 9 0 0 12288 0 1 10 0 0 4
133 353
214 353
214 369
342 369
2 1 10 0 0 4224 0 20 10 0 0 4
254 294
334 294
334 351
342 351
1 2 11 0 0 12288 0 3 11 0 0 4
131 206
193 206
193 314
340 314
2 1 12 0 0 8320 0 22 11 0 0 4
253 153
309 153
309 296
340 296
3 2 13 0 0 4224 0 13 12 0 0 4
479 290
707 290
707 255
715 255
3 1 8 0 0 0 0 16 12 0 0 4
480 163
570 163
570 237
715 237
1 2 9 0 0 12416 0 1 13 0 0 6
133 353
199 353
199 274
416 274
416 299
424 299
1 1 14 0 0 12416 0 2 13 0 0 4
135 302
204 302
204 281
424 281
3 2 15 0 0 12416 0 18 14 0 0 6
375 146
421 146
421 183
709 183
709 165
717 165
3 1 16 0 0 4224 0 15 14 0 0 4
619 162
709 162
709 147
717 147
3 2 17 0 0 4224 0 17 15 0 0 4
374 200
566 200
566 171
574 171
3 1 8 0 0 0 0 16 15 0 0 4
480 163
566 163
566 153
574 153
1 2 11 0 0 12416 0 3 16 0 0 4
131 206
205 206
205 172
425 172
1 1 18 0 0 12416 0 4 16 0 0 6
132 156
203 156
203 168
417 168
417 154
425 154
2 2 19 0 0 8320 0 19 17 0 0 4
254 350
321 350
321 209
329 209
1 1 14 0 0 0 0 2 17 0 0 6
135 302
215 302
215 183
316 183
316 191
329 191
2 2 20 0 0 4224 0 21 18 0 0 4
255 198
322 198
322 155
330 155
1 1 18 0 0 0 0 4 18 0 0 4
132 156
213 156
213 137
330 137
1 1 9 0 0 0 0 1 19 0 0 4
133 353
210 353
210 350
218 350
1 1 14 0 0 0 0 2 20 0 0 4
135 302
210 302
210 294
218 294
1 1 11 0 0 0 0 3 21 0 0 4
131 206
211 206
211 198
219 198
1 1 18 0 0 0 0 4 22 0 0 4
132 156
209 156
209 153
217 153
8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
461 64 610 88
471 72 599 88
16 2 BIT COMPARATOR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
929 317 974 341
939 325 963 341
3 A<B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
933 215 978 239
943 223 967 239
3 A=B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
931 111 976 135
941 119 965 135
3 A>B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
72 336 109 360
82 344 98 360
2 B0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
72 276 109 300
82 284 98 300
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
71 182 108 206
81 190 97 206
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
74 140 111 164
84 148 100 164
2 A1
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
