CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
190 40 5 140 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 599 250 0 1 11
0 2
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 203 258 0 1 11
0 3
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89855e-315 0
0
12 Hex Display~
7 693 82 0 18 19
10 8 9 10 11 0 0 0 0 0
0 0 1 1 0 0 1 1 4
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3124 0 0
2
5.89855e-315 0
0
12 Hex Display~
7 315 86 0 18 19
10 4 5 6 7 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3421 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 516 149 0 3 22
0 13 14 12
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U3C
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
8157 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 317 167 0 3 22
0 5 5 13
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U3B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
5572 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 691 159 0 3 22
0 11 11 14
0
0 0 608 180
6 74LS08
-21 -24 21 -16
3 U3A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
8901 0 0
2
5.89855e-315 0
0
7 Pulser~
4 593 368 0 10 12
0 16 17 15 18 0 0 5 5 5
8
0
0 0 4640 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7361 0 0
2
5.89855e-315 0
0
6 74LS90
107 687 284 0 10 21
0 2 2 12 12 15 8 11 10 9
8
0
0 0 4832 0
6 74LS90
-21 -51 21 -43
2 U2
-7 -52 7 -44
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
4747 0 0
2
5.89855e-315 0
0
6 74LS90
107 315 289 0 10 21
0 3 3 12 12 11 4 7 6 5
4
0
0 0 4832 0
6 74LS90
-21 -51 21 -43
2 U1
-7 -52 7 -44
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
972 0 0
2
5.89855e-315 0
0
26
1 2 2 0 0 4096 0 1 9 0 0 4
611 250
636 250
636 266
655 266
1 1 2 0 0 4224 0 1 9 0 0 4
611 250
641 250
641 257
655 257
1 2 3 0 0 4096 0 2 10 0 0 4
215 258
259 258
259 271
283 271
1 1 3 0 0 4224 0 2 10 0 0 4
215 258
264 258
264 262
283 262
10 1 4 0 0 8320 0 10 4 0 0 5
347 316
386 316
386 138
324 138
324 110
9 2 5 0 0 8320 0 10 4 0 0 5
347 298
381 298
381 133
318 133
318 110
8 3 6 0 0 8320 0 10 4 0 0 5
347 280
376 280
376 123
312 123
312 110
7 4 7 0 0 8320 0 10 4 0 0 5
347 262
371 262
371 118
306 118
306 110
10 1 8 0 0 8320 0 9 3 0 0 5
719 311
753 311
753 129
702 129
702 106
9 2 9 0 0 8320 0 9 3 0 0 5
719 293
748 293
748 124
696 124
696 106
8 3 10 0 0 8320 0 9 3 0 0 5
719 275
743 275
743 119
690 119
690 106
7 4 11 0 0 8192 0 9 3 0 0 5
719 257
738 257
738 114
684 114
684 106
3 4 12 0 0 12288 0 5 9 0 0 4
489 149
482 149
482 284
655 284
3 3 12 0 0 0 0 5 9 0 0 4
489 149
487 149
487 275
655 275
3 4 12 0 0 8320 0 5 10 0 0 6
489 149
366 149
366 341
259 341
259 289
283 289
3 3 12 0 0 0 0 5 10 0 0 6
489 149
361 149
361 242
269 242
269 280
283 280
3 1 13 0 0 12416 0 6 5 0 0 6
290 167
288 167
288 129
549 129
549 158
534 158
3 2 14 0 0 4224 0 7 5 0 0 4
664 159
544 159
544 140
534 140
9 2 5 0 0 0 0 10 6 0 0 4
347 298
356 298
356 158
335 158
9 1 5 0 0 0 0 10 6 0 0 4
347 298
351 298
351 176
335 176
7 2 11 0 0 0 0 9 7 0 0 4
719 257
733 257
733 150
709 150
7 1 11 0 0 0 0 9 7 0 0 4
719 257
723 257
723 168
709 168
10 6 4 0 0 0 0 10 10 0 0 6
347 316
351 316
351 336
264 336
264 316
277 316
7 5 11 0 0 12416 0 9 10 0 0 6
719 257
728 257
728 331
269 331
269 307
277 307
10 6 8 0 0 0 0 9 9 0 0 6
719 311
723 311
723 326
636 326
636 311
649 311
3 5 15 0 0 8320 0 8 9 0 0 4
617 359
641 359
641 302
649 302
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
396 417 577 441
406 425 566 441
20 DIVIDE BY 27 COUNTER
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
