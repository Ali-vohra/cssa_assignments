CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
350 120 4 220 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
4
13 Logic Switch~
5 362 233 0 1 11
0 6
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89855e-315 0
0
12 Hex Display~
7 632 158 0 18 19
10 2 3 4 5 0 0 0 0 0
0 1 1 1 0 0 0 0 7
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
391 0 0
2
5.89855e-315 0
0
7 Pulser~
4 384 332 0 10 12
0 8 9 7 10 0 0 5 5 1
8
0
0 0 4640 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3124 0 0
2
5.89855e-315 0
0
6 74LS90
107 494 260 0 10 21
0 6 6 6 6 7 2 5 4 3
2
0
0 0 4832 0
6 74LS90
-21 -51 21 -43
2 U1
-7 -52 7 -44
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
3421 0 0
2
5.89855e-315 0
0
10
10 1 2 0 0 4224 0 4 2 0 0 3
526 287
641 287
641 182
9 2 3 0 0 4224 0 4 2 0 0 3
526 269
635 269
635 182
8 3 4 0 0 4224 0 4 2 0 0 3
526 251
629 251
629 182
7 4 5 0 0 4224 0 4 2 0 0 3
526 233
623 233
623 182
1 4 6 0 0 4096 0 1 4 0 0 4
374 233
438 233
438 260
462 260
1 3 6 0 0 4096 0 1 4 0 0 4
374 233
443 233
443 251
462 251
1 2 6 0 0 4096 0 1 4 0 0 4
374 233
448 233
448 242
462 242
1 1 6 0 0 4224 0 1 4 0 0 2
374 233
462 233
10 6 2 0 0 0 0 4 4 0 0 6
526 287
530 287
530 302
443 302
443 287
456 287
3 5 7 0 0 8320 0 3 4 0 0 4
408 323
448 323
448 278
456 278
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 19
432 361 612 385
436 364 607 380
19 DIVIDE BY 9 COUNTER
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
