CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
40 10 30 70 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 E:\CM60S\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
143654930 0
0
6 Title:
5 Name:
0
0
0
38
13 Logic Switch~
5 331 124 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V11
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
43331.8 0
0
13 Logic Switch~
5 494 234 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V10
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
43331.8 1
0
13 Logic Switch~
5 592 93 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
43331.8 2
0
13 Logic Switch~
5 89 531 0 10 11
0 35 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
43331.8 3
0
13 Logic Switch~
5 91 479 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8157 0 0
2
43331.8 4
0
13 Logic Switch~
5 90 430 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5572 0 0
2
43331.8 5
0
13 Logic Switch~
5 92 381 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8901 0 0
2
43331.8 6
0
13 Logic Switch~
5 98 257 0 10 11
0 31 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7361 0 0
2
43331.8 7
0
13 Logic Switch~
5 97 204 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4747 0 0
2
43331.8 8
0
13 Logic Switch~
5 96 152 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
972 0 0
2
43331.8 9
0
13 Logic Switch~
5 96 104 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3472 0 0
2
43331.8 10
0
14 Logic Display~
6 964 173 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9998 0 0
2
43331.8 11
0
14 Logic Display~
6 965 233 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3536 0 0
2
43331.8 12
0
9 2-In AND~
219 221 804 0 3 22
0 11 10 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
4597 0 0
2
43331.8 13
0
14 Logic Display~
6 967 281 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3835 0 0
2
43331.8 14
0
9 2-In AND~
219 221 761 0 3 22
0 15 10 13
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
3670 0 0
2
43331.8 15
0
9 2-In AND~
219 220 702 0 3 22
0 11 17 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
5616 0 0
2
43331.8 16
0
14 Logic Display~
6 967 331 0 1 2
10 19
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9323 0 0
2
43331.8 17
0
9 2-In AND~
219 219 651 0 3 22
0 10 23 22
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
317 0 0
2
43331.8 18
0
9 2-In AND~
219 219 599 0 3 22
0 15 17 24
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
3108 0 0
2
43331.8 19
0
9 2-In AND~
219 219 551 0 3 22
0 11 26 25
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
4299 0 0
2
43331.8 20
0
14 Logic Display~
6 965 382 0 1 2
10 27
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9672 0 0
2
43331.8 21
0
6 74LS83
105 708 96 0 14 29
0 9 14 20 29 8 13 4 28 4
7 12 19 27 6
0
0 0 13040 0
7 74LS83A
-24 -60 25 -52
2 U6
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
7876 0 0
2
43331.8 22
0
9 2-In AND~
219 219 503 0 3 22
0 10 31 30
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
6369 0 0
2
43331.8 23
0
9 2-In AND~
219 218 456 0 3 22
0 23 17 32
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
9172 0 0
2
43331.8 24
0
9 2-In AND~
219 217 406 0 3 22
0 15 26 33
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
7100 0 0
2
43331.8 25
0
9 2-In AND~
219 217 358 0 3 22
0 11 35 34
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
3820 0 0
2
43331.8 26
0
14 Logic Display~
6 967 428 0 1 2
10 36
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7678 0 0
2
43331.8 27
0
6 74LS83
105 595 229 0 14 29
0 18 21 32 38 16 22 30 37 3
14 20 28 36 9
0
0 0 13040 0
7 74LS83A
-24 -60 25 -52
2 U4
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
961 0 0
2
43331.8 28
0
9 2-In AND~
219 216 304 0 3 22
0 31 17 37
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3178 0 0
2
43331.8 29
0
14 Logic Display~
6 968 476 0 1 2
10 39
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3409 0 0
2
43331.8 30
0
9 2-In AND~
219 215 254 0 3 22
0 23 26 40
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3951 0 0
2
43331.8 31
0
9 2-In AND~
219 216 202 0 3 22
0 15 35 41
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
8885 0 0
2
43331.8 32
0
9 2-In AND~
219 216 149 0 3 22
0 31 26 42
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3780 0 0
2
43331.8 33
0
9 2-In AND~
219 216 95 0 3 22
0 23 35 43
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
9265 0 0
2
43331.8 34
0
6 74LS83
105 455 133 0 14 29
0 25 34 41 43 24 33 40 42 2
21 29 38 39 18
0
0 0 13040 0
7 74LS83A
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
9442 0 0
2
43331.8 35
0
14 Logic Display~
6 966 532 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9424 0 0
2
43331.8 36
0
9 2-In AND~
219 216 41 0 3 22
0 31 35 5
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
9968 0 0
2
43331.8 37
0
67
1 9 2 0 0 4224 0 1 36 0 0 4
343 124
415 124
415 178
423 178
1 9 3 0 0 4224 0 2 29 0 0 4
506 234
555 234
555 274
563 274
1 9 4 0 0 4224 0 3 23 0 0 4
604 93
668 93
668 141
676 141
3 1 5 0 0 4224 0 38 37 0 0 7
237 41
905 41
905 517
882 517
882 558
966 558
966 550
14 1 6 0 0 4224 0 23 12 0 0 5
740 141
877 141
877 203
964 203
964 191
10 1 7 0 0 8320 0 23 13 0 0 5
740 87
877 87
877 255
965 255
965 251
3 5 8 0 0 8320 0 14 23 0 0 4
242 804
668 804
668 96
676 96
14 1 9 0 0 8320 0 29 23 0 0 4
627 274
668 274
668 60
676 60
1 2 10 0 0 8320 0 7 14 0 0 4
104 381
189 381
189 813
197 813
1 1 11 0 0 8320 0 11 14 0 0 4
108 104
187 104
187 795
197 795
11 1 12 0 0 8320 0 23 15 0 0 5
740 96
877 96
877 305
967 305
967 299
3 6 13 0 0 8320 0 16 23 0 0 4
242 761
668 761
668 105
676 105
10 2 14 0 0 8320 0 29 23 0 0 4
627 220
668 220
668 69
676 69
1 2 10 0 0 0 0 7 16 0 0 4
104 381
189 381
189 770
197 770
1 1 15 0 0 8320 0 10 16 0 0 4
108 152
187 152
187 752
197 752
3 5 16 0 0 8320 0 17 29 0 0 4
241 702
555 702
555 229
563 229
1 1 11 0 0 0 0 11 17 0 0 4
108 104
186 104
186 693
196 693
1 2 17 0 0 8320 0 6 17 0 0 4
102 430
188 430
188 711
196 711
14 1 18 0 0 4224 0 36 29 0 0 4
487 178
555 178
555 193
563 193
12 1 19 0 0 8320 0 23 18 0 0 5
740 105
878 105
878 357
967 357
967 349
1 7 4 0 0 0 0 3 23 0 0 4
604 93
668 93
668 114
676 114
11 3 20 0 0 8320 0 29 23 0 0 4
627 229
668 229
668 78
676 78
10 2 21 0 0 8320 0 36 29 0 0 4
487 124
555 124
555 202
563 202
3 6 22 0 0 8320 0 19 29 0 0 4
240 651
555 651
555 238
563 238
1 2 23 0 0 8320 0 9 19 0 0 4
109 204
187 204
187 660
195 660
1 1 10 0 0 0 0 7 19 0 0 4
104 381
187 381
187 642
195 642
3 5 24 0 0 8320 0 20 36 0 0 4
240 599
415 599
415 133
423 133
1 2 17 0 0 0 0 6 20 0 0 4
102 430
187 430
187 608
195 608
1 1 15 0 0 0 0 10 20 0 0 4
108 152
187 152
187 590
195 590
3 1 25 0 0 8320 0 21 36 0 0 4
240 551
415 551
415 97
423 97
1 2 26 0 0 4096 0 5 21 0 0 4
103 479
187 479
187 560
195 560
1 1 11 0 0 0 0 11 21 0 0 4
108 104
187 104
187 542
195 542
13 1 27 0 0 8320 0 23 22 0 0 5
740 114
878 114
878 407
965 407
965 400
12 8 28 0 0 8320 0 29 23 0 0 4
627 238
668 238
668 123
676 123
11 4 29 0 0 4224 0 36 23 0 0 4
487 133
668 133
668 87
676 87
3 7 30 0 0 4224 0 24 29 0 0 4
240 503
555 503
555 247
563 247
1 2 31 0 0 8320 0 8 24 0 0 4
110 257
187 257
187 512
195 512
1 1 10 0 0 0 0 7 24 0 0 4
104 381
187 381
187 494
195 494
3 3 32 0 0 4224 0 25 29 0 0 4
239 456
555 456
555 211
563 211
1 2 17 0 0 0 0 6 25 0 0 4
102 430
186 430
186 465
194 465
1 1 23 0 0 0 0 9 25 0 0 4
109 204
186 204
186 447
194 447
3 6 33 0 0 8320 0 26 36 0 0 4
238 406
415 406
415 142
423 142
1 2 26 0 0 0 0 5 26 0 0 4
103 479
185 479
185 415
193 415
1 1 15 0 0 0 0 10 26 0 0 4
108 152
185 152
185 397
193 397
3 2 34 0 0 8320 0 27 36 0 0 4
238 358
415 358
415 106
423 106
1 2 35 0 0 8192 0 4 27 0 0 4
101 531
185 531
185 367
193 367
1 1 11 0 0 0 0 11 27 0 0 4
108 104
185 104
185 349
193 349
13 1 36 0 0 4224 0 29 28 0 0 5
627 247
879 247
879 457
967 457
967 446
3 8 37 0 0 4224 0 30 29 0 0 4
237 304
555 304
555 256
563 256
12 4 38 0 0 8320 0 36 29 0 0 4
487 142
555 142
555 220
563 220
1 2 17 0 0 0 0 6 30 0 0 4
102 430
184 430
184 313
192 313
1 1 31 0 0 0 0 8 30 0 0 4
110 257
184 257
184 295
192 295
13 1 39 0 0 4224 0 36 31 0 0 5
487 151
880 151
880 507
968 507
968 494
3 7 40 0 0 4224 0 32 36 0 0 4
236 254
415 254
415 151
423 151
1 2 26 0 0 8192 0 5 32 0 0 4
103 479
183 479
183 263
191 263
1 1 23 0 0 0 0 9 32 0 0 4
109 204
183 204
183 245
191 245
3 3 41 0 0 4224 0 33 36 0 0 4
237 202
415 202
415 115
423 115
1 2 35 0 0 8192 0 4 33 0 0 4
101 531
184 531
184 211
192 211
1 1 15 0 0 0 0 10 33 0 0 4
108 152
184 152
184 193
192 193
3 8 42 0 0 4224 0 34 36 0 0 4
237 149
415 149
415 160
423 160
3 4 43 0 0 4224 0 35 36 0 0 4
237 95
415 95
415 124
423 124
1 2 26 0 0 8320 0 5 34 0 0 4
103 479
184 479
184 158
192 158
1 1 31 0 0 0 0 8 34 0 0 4
110 257
184 257
184 140
192 140
1 2 35 0 0 8192 0 4 35 0 0 4
101 531
184 531
184 104
192 104
1 1 23 0 0 0 0 9 35 0 0 4
109 204
184 204
184 86
192 86
1 2 35 0 0 8320 0 4 38 0 0 4
101 531
184 531
184 50
192 50
1 1 31 0 0 0 0 8 38 0 0 4
110 257
184 257
184 32
192 32
17
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
621 838 763 853
636 850 747 861
16 4 BIT MULTIPLIER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
49 82 73 106
59 90 75 106
2 A3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
49 134 73 158
59 142 75 158
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
50 183 74 207
60 191 76 207
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
49 231 73 255
59 239 75 255
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
46 355 70 379
56 363 72 379
2 B3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
45 405 69 429
55 413 71 429
2 B2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
43 457 67 481
53 465 69 481
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
44 508 68 532
54 516 70 532
2 B0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
976 520 1000 544
986 528 1002 544
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
976 464 1000 488
986 472 1002 488
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
977 417 1001 441
987 425 1003 441
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
976 363 1000 387
986 371 1002 387
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
976 321 1000 345
986 329 1002 345
2 S4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
973 220 993 235
987 232 1001 243
2 S6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
975 160 995 175
989 171 1003 182
2 S7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
980 272 1004 296
985 276 1001 292
2 S5
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
