CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 10 30 70 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
24
13 Logic Switch~
5 329 586 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V5
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3409 0 0
2
43362 0
0
13 Logic Switch~
5 279 587 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V4
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3951 0 0
2
43362 0
0
13 Logic Switch~
5 224 586 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V3
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8885 0 0
2
43362 0
0
13 Logic Switch~
5 156 587 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V2
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3780 0 0
2
43362 0
0
13 Logic Switch~
5 118 252 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9265 0 0
2
43362 0
0
9 Inverter~
13 133 516 0 2 22
0 2 3
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U3A
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
9442 0 0
2
43362 0
0
14 Logic Display~
6 753 812 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L16
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9424 0 0
2
43362 0
0
14 Logic Display~
6 757 765 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L15
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9968 0 0
2
43362 0
0
14 Logic Display~
6 756 713 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L14
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9281 0 0
2
43362 0
0
14 Logic Display~
6 756 666 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L13
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8464 0 0
2
43362 0
0
14 Logic Display~
6 758 617 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7168 0 0
2
43362 0
0
14 Logic Display~
6 759 562 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3171 0 0
2
43362 0
0
14 Logic Display~
6 759 511 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4139 0 0
2
43362 0
0
14 Logic Display~
6 762 457 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6435 0 0
2
43362 0
0
14 Logic Display~
6 761 402 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5283 0 0
2
43362 0
0
14 Logic Display~
6 761 347 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6874 0 0
2
43362 0
0
14 Logic Display~
6 761 292 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5305 0 0
2
43362 0
0
14 Logic Display~
6 760 242 0 1 2
10 18
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
34 0 0
2
43362 0
0
14 Logic Display~
6 759 186 0 1 2
10 19
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
969 0 0
2
43362 0
0
14 Logic Display~
6 757 131 0 1 2
10 20
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8402 0 0
2
43362 0
0
14 Logic Display~
6 757 81 0 1 2
10 21
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3751 0 0
2
43362 0
0
14 Logic Display~
6 756 32 0 1 2
10 22
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4292 0 0
2
43362 0
0
10 1x8 DEMUX~
94 377 116 0 13 27
0 2 23 6 5 4 22 21 20 19
18 17 16 15
9 1x8 DEMUX
1 0 528 0
0
2 U1
1 -68 15 -60
0
0
0
0
0
0
27

0 1 4 6 7 8 9 10 11 12
13 14 15 16 1 4 6 7 8 9
10 11 12 13 14 15 16 0
0 0 0 0 0 0 0 0
1 U
6118 0 0
2
43362 0
0
10 1x8 DEMUX~
94 375 392 0 13 27
0 3 23 6 5 4 14 13 12 11
10 9 8 7
9 1x8 DEMUX
2 0 528 0
0
2 U2
1 -68 15 -60
0
0
0
0
0
0
27

0 1 4 6 7 8 9 10 11 12
13 14 15 16 1 4 6 7 8 9
10 11 12 13 14 15 16 0
0 0 0 0 0 0 0 0
1 U
34 0 0
2
43362 0
0
27
1 1 2 0 0 4224 0 4 23 0 0 3
157 574
157 81
344 81
2 1 3 0 0 8320 0 6 24 0 0 3
136 498
136 357
342 357
1 1 2 0 0 0 0 6 4 0 0 4
136 534
136 567
157 567
157 574
1 5 4 0 0 4096 0 1 24 0 0 3
330 573
330 438
342 438
1 4 5 0 0 4096 0 2 24 0 0 3
280 574
280 427
342 427
1 3 6 0 0 4096 0 3 24 0 0 3
225 573
225 415
342 415
1 5 4 0 0 4224 0 1 23 0 0 3
330 573
330 162
344 162
1 4 5 0 0 4224 0 2 23 0 0 3
280 574
280 151
344 151
1 3 6 0 0 4224 0 3 23 0 0 3
225 573
225 139
344 139
13 1 7 0 0 8320 0 24 7 0 0 4
424 357
563 357
563 830
753 830
12 1 8 0 0 8320 0 24 8 0 0 4
424 369
576 369
576 783
757 783
11 1 9 0 0 8320 0 24 9 0 0 4
424 381
589 381
589 731
756 731
10 1 10 0 0 8320 0 24 10 0 0 4
424 392
600 392
600 684
756 684
9 1 11 0 0 8320 0 24 11 0 0 4
424 403
613 403
613 635
758 635
8 1 12 0 0 4224 0 24 12 0 0 4
424 415
626 415
626 580
759 580
7 1 13 0 0 4224 0 24 13 0 0 4
424 427
636 427
636 529
759 529
6 1 14 0 0 4224 0 24 14 0 0 5
424 438
709 438
709 484
762 484
762 475
13 1 15 0 0 8320 0 23 15 0 0 4
426 81
644 81
644 420
761 420
12 1 16 0 0 8320 0 23 16 0 0 4
426 93
656 93
656 365
761 365
11 1 17 0 0 4224 0 23 17 0 0 4
426 105
667 105
667 310
761 310
10 1 18 0 0 4224 0 23 18 0 0 4
426 116
680 116
680 260
760 260
9 1 19 0 0 4224 0 23 19 0 0 5
426 127
689 127
689 214
759 214
759 204
8 1 20 0 0 4224 0 23 20 0 0 5
426 139
694 139
694 159
757 159
757 149
7 1 21 0 0 4224 0 23 21 0 0 5
426 151
699 151
699 106
757 106
757 99
6 1 22 0 0 4224 0 23 22 0 0 5
426 162
703 162
703 58
756 58
756 50
1 2 23 0 0 4096 0 5 24 0 0 4
130 252
329 252
329 392
342 392
1 2 23 0 0 4224 0 5 23 0 0 4
130 252
336 252
336 116
344 116
21
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
775 793 820 808
790 804 804 815
2 D0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
779 749 822 764
793 761 807 772
2 D1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
780 695 825 710
795 707 809 718
2 D2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
780 649 823 664
794 660 808 671
2 D3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
781 598 824 613
795 609 809 620
2 D4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
783 544 826 559
797 556 811 567
2 D5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
785 493 828 508
799 505 813 516
2 D6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
786 439 829 454
800 451 814 462
2 D7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
788 386 833 401
803 397 817 408
2 D8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
787 329 830 344
801 340 815 351
2 D9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
789 277 839 292
803 289 824 300
3 D10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
790 224 840 239
804 236 825 247
3 D11
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
790 170 840 185
804 181 825 192
3 D12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
791 117 841 132
805 129 826 140
3 D13
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
790 67 842 82
805 79 826 90
3 D14
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
791 14 841 29
805 26 826 37
3 D15
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
310 607 353 622
324 618 338 629
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
257 606 300 621
271 617 285 628
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
203 607 246 622
217 618 231 629
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
134 607 179 622
149 618 163 629
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
66 230 102 245
80 242 87 253
1 A
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
