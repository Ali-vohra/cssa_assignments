CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 300 30 110 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
24
13 Logic Switch~
5 703 223 0 1 11
0 7
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 382 378 0 1 11
0 18
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 115 245 0 10 11
0 35 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3124 0 0
2
5.89855e-315 0
0
13 Logic Switch~
5 86 450 0 1 11
0 19
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.89855e-315 0
0
14 Logic Display~
6 977 328 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8157 0 0
2
5.89855e-315 0
0
12 Hex Display~
7 1025 91 0 16 19
10 3 4 5 6 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
5572 0 0
2
5.89855e-315 0
0
9 Inverter~
13 556 481 0 2 22
0 9 8
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
8901 0 0
2
5.89855e-315 0
0
5 4030~
219 728 517 0 3 22
0 14 8 10
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U8D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 4 0
1 U
7361 0 0
2
5.89855e-315 0
0
5 4030~
219 728 466 0 3 22
0 15 8 11
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U8C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 4 0
1 U
4747 0 0
2
5.89855e-315 0
0
5 4030~
219 728 411 0 3 22
0 16 8 12
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U8B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 4 0
1 U
972 0 0
2
5.89855e-315 0
0
5 4030~
219 727 358 0 3 22
0 17 8 13
0
0 0 608 0
4 4030
-7 -24 21 -16
3 U8A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
3472 0 0
2
5.89855e-315 0
0
6 74LS83
105 845 284 0 14 29
0 8 7 8 7 13 12 11 10 9
6 5 4 3 2
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U7
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
9998 0 0
2
5.89855e-315 0
0
8 3-In OR~
219 491 412 0 4 22
0 21 20 22 9
0
0 0 608 270
4 4075
-14 -24 14 -16
3 U6A
28 -7 49 1
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 3 0
1 U
3536 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 535 357 0 3 22
0 23 24 21
0
0 0 608 270
6 74LS08
-21 -24 21 -16
3 U5B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
4597 0 0
2
5.89855e-315 0
0
9 2-In AND~
219 455 358 0 3 22
0 25 24 22
0
0 0 608 270
6 74LS08
-21 -24 21 -16
3 U5A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3835 0 0
2
5.89855e-315 0
0
6 74LS83
105 627 288 0 14 29
0 24 25 23 26 18 9 9 18 18
17 16 15 14 44
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U4
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
3670 0 0
2
5.89855e-315 0
0
8 Hex Key~
166 290 95 0 11 12
0 27 28 29 30 0 0 0 0 0
9 57
0
0 0 4640 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
5616 0 0
2
5.89855e-315 0
0
6 74LS83
105 380 289 0 14 29
0 30 29 28 27 34 33 32 31 19
24 25 23 26 20
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U3
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
9323 0 0
2
5.89855e-315 0
0
8 Hex Key~
166 59 99 0 11 12
0 37 39 41 43 0 0 0 0 0
9 57
0
0 0 4640 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
317 0 0
2
5.89855e-315 0
0
9 Inverter~
13 86 409 0 2 22
0 37 36
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
3108 0 0
2
5.89855e-315 0
0
9 Inverter~
13 86 369 0 2 22
0 39 38
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
4299 0 0
2
5.89855e-315 0
0
9 Inverter~
13 86 329 0 2 22
0 41 40
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
9672 0 0
2
5.89855e-315 0
0
9 Inverter~
13 85 288 0 2 22
0 43 42
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
7876 0 0
2
5.89855e-315 0
0
6 74LS83
105 210 290 0 14 29
0 35 19 35 19 42 40 38 36 19
34 33 32 31 45
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
6369 0 0
2
5.89855e-315 0
0
61
14 1 2 0 0 4224 0 12 5 0 0 5
877 329
965 329
965 354
977 354
977 346
13 1 3 0 0 8320 0 12 6 0 0 3
877 302
1034 302
1034 115
12 2 4 0 0 8320 0 12 6 0 0 3
877 293
1028 293
1028 115
11 3 5 0 0 8320 0 12 6 0 0 3
877 284
1022 284
1022 115
10 4 6 0 0 8320 0 12 6 0 0 3
877 275
1016 275
1016 115
1 4 7 0 0 4096 0 1 12 0 0 4
715 223
800 223
800 275
813 275
1 2 7 0 0 4224 0 1 12 0 0 4
715 223
805 223
805 257
813 257
2 3 8 0 0 8192 0 7 12 0 0 4
577 481
681 481
681 266
813 266
2 1 8 0 0 8320 0 7 12 0 0 4
577 481
706 481
706 248
813 248
4 9 9 0 0 8320 0 13 12 0 0 5
494 442
494 444
785 444
785 329
813 329
3 8 10 0 0 8320 0 8 12 0 0 4
761 517
790 517
790 311
813 311
3 7 11 0 0 8320 0 9 12 0 0 4
761 466
795 466
795 302
813 302
3 6 12 0 0 8320 0 10 12 0 0 4
761 411
800 411
800 293
813 293
3 5 13 0 0 8320 0 11 12 0 0 4
760 358
805 358
805 284
813 284
2 2 8 0 0 0 0 7 8 0 0 4
577 481
684 481
684 526
712 526
2 2 8 0 0 0 0 7 9 0 0 4
577 481
694 481
694 475
712 475
2 2 8 0 0 0 0 7 10 0 0 4
577 481
699 481
699 420
712 420
2 2 8 0 0 0 0 7 11 0 0 4
577 481
703 481
703 367
711 367
4 1 9 0 0 0 0 13 7 0 0 3
494 442
494 481
541 481
13 1 14 0 0 8320 0 16 8 0 0 4
659 306
689 306
689 508
712 508
12 1 15 0 0 8320 0 16 9 0 0 4
659 297
694 297
694 457
712 457
11 1 16 0 0 8320 0 16 10 0 0 4
659 288
699 288
699 402
712 402
10 1 17 0 0 8320 0 16 11 0 0 4
659 279
703 279
703 349
711 349
1 9 18 0 0 12288 0 2 16 0 0 6
394 378
424 378
424 331
577 331
577 333
595 333
1 8 18 0 0 12416 0 2 16 0 0 4
394 378
429 378
429 315
595 315
1 5 18 0 0 0 0 2 16 0 0 4
394 378
434 378
434 288
595 288
1 9 19 0 0 4224 0 4 18 0 0 4
98 450
340 450
340 334
348 334
4 7 9 0 0 0 0 13 16 0 0 5
494 442
494 444
582 444
582 306
595 306
4 6 9 0 0 0 0 13 16 0 0 5
494 442
494 439
587 439
587 297
595 297
14 2 20 0 0 4224 0 18 13 0 0 3
412 334
494 334
494 397
3 1 21 0 0 8320 0 14 13 0 0 4
533 380
533 384
503 384
503 396
3 3 22 0 0 8320 0 15 13 0 0 4
453 381
453 385
485 385
485 396
12 1 23 0 0 4096 0 18 14 0 0 3
412 298
542 298
542 335
10 2 24 0 0 4096 0 18 14 0 0 3
412 280
524 280
524 335
11 1 25 0 0 4096 0 18 15 0 0 3
412 289
462 289
462 336
10 2 24 0 0 0 0 18 15 0 0 3
412 280
444 280
444 336
13 4 26 0 0 4224 0 18 16 0 0 4
412 307
572 307
572 279
595 279
12 3 23 0 0 4224 0 18 16 0 0 4
412 298
577 298
577 270
595 270
11 2 25 0 0 4224 0 18 16 0 0 4
412 289
582 289
582 261
595 261
10 1 24 0 0 4224 0 18 16 0 0 4
412 280
587 280
587 252
595 252
1 4 27 0 0 4224 0 17 18 0 0 3
299 119
299 280
348 280
2 3 28 0 0 4224 0 17 18 0 0 3
293 119
293 271
348 271
3 2 29 0 0 4224 0 17 18 0 0 3
287 119
287 262
348 262
4 1 30 0 0 4224 0 17 18 0 0 3
281 119
281 253
348 253
13 8 31 0 0 4224 0 24 18 0 0 4
242 308
340 308
340 316
348 316
12 7 32 0 0 4224 0 24 18 0 0 4
242 299
340 299
340 307
348 307
11 6 33 0 0 4224 0 24 18 0 0 4
242 290
340 290
340 298
348 298
10 5 34 0 0 4224 0 24 18 0 0 4
242 281
340 281
340 289
348 289
1 4 19 0 0 0 0 4 24 0 0 4
98 450
150 450
150 281
178 281
1 2 19 0 0 0 0 4 24 0 0 4
98 450
155 450
155 263
178 263
1 3 35 0 0 4096 0 3 24 0 0 4
127 245
165 245
165 272
178 272
1 1 35 0 0 4224 0 3 24 0 0 4
127 245
170 245
170 254
178 254
1 9 19 0 0 0 0 4 24 0 0 4
98 450
170 450
170 335
178 335
2 8 36 0 0 8320 0 20 24 0 0 4
107 409
160 409
160 317
178 317
1 1 37 0 0 4224 0 19 20 0 0 5
68 123
68 274
53 274
53 409
71 409
2 7 38 0 0 8320 0 21 24 0 0 4
107 369
165 369
165 308
178 308
2 1 39 0 0 4224 0 19 21 0 0 3
62 123
62 369
71 369
2 6 40 0 0 4224 0 22 24 0 0 4
107 329
170 329
170 299
178 299
3 1 41 0 0 4224 0 19 22 0 0 3
56 123
56 329
71 329
2 5 42 0 0 4224 0 23 24 0 0 4
106 288
170 288
170 290
178 290
4 1 43 0 0 4224 0 19 23 0 0 3
50 123
50 288
70 288
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
428 570 607 592
437 577 597 593
20 BCD SUBTRACTOR (9'S)
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
